// av_sata_xcvr_core.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module av_sata_xcvr_core (
		input  wire [0:0]  pll_powerdown,           //           pll_powerdown.pll_powerdown
		input  wire [0:0]  tx_analogreset,          //          tx_analogreset.tx_analogreset
		input  wire [0:0]  tx_digitalreset,         //         tx_digitalreset.tx_digitalreset
		output wire [0:0]  tx_serial_data,          //          tx_serial_data.tx_serial_data
		input  wire [0:0]  ext_pll_clk,             //             ext_pll_clk.ext_pll_clk
		input  wire [0:0]  rx_analogreset,          //          rx_analogreset.rx_analogreset
		input  wire [0:0]  rx_digitalreset,         //         rx_digitalreset.rx_digitalreset
		input  wire [0:0]  rx_cdr_refclk,           //           rx_cdr_refclk.rx_cdr_refclk
		input  wire [0:0]  rx_serial_data,          //          rx_serial_data.rx_serial_data
		output wire [0:0]  rx_is_lockedtoref,       //       rx_is_lockedtoref.rx_is_lockedtoref
		output wire [0:0]  rx_is_lockedtodata,      //      rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [0:0]  tx_std_coreclkin,        //        tx_std_coreclkin.tx_std_coreclkin
		input  wire [0:0]  rx_std_coreclkin,        //        rx_std_coreclkin.rx_std_coreclkin
		output wire [0:0]  tx_std_clkout,           //           tx_std_clkout.tx_std_clkout
		output wire [0:0]  rx_std_clkout,           //           rx_std_clkout.rx_std_clkout
		input  wire [0:0]  tx_std_elecidle,         //         tx_std_elecidle.tx_std_elecidle
		output wire [0:0]  rx_std_signaldetect,     //     rx_std_signaldetect.rx_std_signaldetect
		output wire [0:0]  tx_cal_busy,             //             tx_cal_busy.tx_cal_busy
		output wire [0:0]  rx_cal_busy,             //             rx_cal_busy.rx_cal_busy
		input  wire [69:0] reconfig_to_xcvr,        //        reconfig_to_xcvr.reconfig_to_xcvr
		output wire [45:0] reconfig_from_xcvr,      //      reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [31:0] tx_parallel_data,        //        tx_parallel_data.tx_parallel_data
		input  wire [3:0]  tx_datak,                //                tx_datak.tx_datak
		input  wire [7:0]  unused_tx_parallel_data, // unused_tx_parallel_data.unused_tx_parallel_data
		output wire [31:0] rx_parallel_data,        //        rx_parallel_data.rx_parallel_data
		output wire [3:0]  rx_datak,                //                rx_datak.rx_datak
		output wire [3:0]  rx_errdetect,            //            rx_errdetect.rx_errdetect
		output wire [3:0]  rx_disperr,              //              rx_disperr.rx_disperr
		output wire [3:0]  rx_runningdisp,          //          rx_runningdisp.rx_runningdisp
		output wire [3:0]  rx_patterndetect,        //        rx_patterndetect.rx_patterndetect
		output wire [3:0]  rx_syncstatus,           //           rx_syncstatus.rx_syncstatus
		output wire [7:0]  unused_rx_parallel_data  // unused_rx_parallel_data.unused_rx_parallel_data
	);

	wire  [63:0] av_sata_xcvr_core_inst_rx_parallel_data; // port fragment

	altera_xcvr_native_av #(
		.tx_enable                       (1),
		.rx_enable                       (1),
		.enable_std                      (1),
		.data_path_select                ("standard"),
		.channels                        (1),
		.bonded_mode                     ("non_bonded"),
		.data_rate                       ("1500 Mbps"),
		.pma_width                       (20),
		.tx_pma_clk_div                  (4),
		.pll_reconfig_enable             (0),
		.pll_external_enable             (1),
		.pll_data_rate                   ("6000 Mbps"),
		.pll_type                        ("CMU"),
		.pma_bonding_mode                ("x1"),
		.plls                            (1),
		.pll_select                      (0),
		.pll_refclk_cnt                  (1),
		.pll_refclk_select               ("0"),
		.pll_refclk_freq                 ("125.0 MHz"),
		.pll_feedback_path               ("internal"),
		.cdr_reconfig_enable             (0),
		.cdr_refclk_cnt                  (1),
		.cdr_refclk_select               (0),
		.cdr_refclk_freq                 ("150.0 MHz"),
		.rx_ppm_detect_threshold         ("1000"),
		.rx_clkslip_enable               (0),
		.std_protocol_hint               ("basic"),
		.std_pcs_pma_width               (20),
		.std_low_latency_bypass_enable   (0),
		.std_tx_pcfifo_mode              ("low_latency"),
		.std_rx_pcfifo_mode              ("low_latency"),
		.std_rx_byte_order_enable        (0),
		.std_rx_byte_order_mode          ("manual"),
		.std_rx_byte_order_width         (9),
		.std_rx_byte_order_symbol_count  (1),
		.std_rx_byte_order_pattern       ("0"),
		.std_rx_byte_order_pad           ("0"),
		.std_tx_byte_ser_enable          (1),
		.std_rx_byte_deser_enable        (1),
		.std_tx_8b10b_enable             (1),
		.std_tx_8b10b_disp_ctrl_enable   (0),
		.std_rx_8b10b_enable             (1),
		.std_rx_rmfifo_enable            (0),
		.std_rx_rmfifo_pattern_p         ("00000"),
		.std_rx_rmfifo_pattern_n         ("00000"),
		.std_tx_bitslip_enable           (0),
		.std_rx_word_aligner_mode        ("manual"),
		.std_rx_word_aligner_pattern_len (10),
		.std_rx_word_aligner_pattern     ("17c"),
		.std_rx_word_aligner_rknumber    (3),
		.std_rx_word_aligner_renumber    (3),
		.std_rx_word_aligner_rgnumber    (3),
		.std_rx_run_length_val           (31),
		.std_tx_bitrev_enable            (0),
		.std_rx_bitrev_enable            (0),
		.std_tx_byterev_enable           (0),
		.std_rx_byterev_enable           (0),
		.std_tx_polinv_enable            (0),
		.std_rx_polinv_enable            (0)
	) av_sata_xcvr_core_inst (
		.pll_powerdown             (pll_powerdown),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       pll_powerdown.pll_powerdown
		.tx_analogreset            (tx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     tx_digitalreset.tx_digitalreset
		.tx_serial_data            (tx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      tx_serial_data.tx_serial_data
		.ext_pll_clk               (ext_pll_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         ext_pll_clk.ext_pll_clk
		.rx_analogreset            (rx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      rx_analogreset.rx_analogreset
		.rx_digitalreset           (rx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     rx_digitalreset.rx_digitalreset
		.rx_cdr_refclk             (rx_cdr_refclk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       rx_cdr_refclk.rx_cdr_refclk
		.rx_serial_data            (rx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      rx_serial_data.rx_serial_data
		.rx_is_lockedtoref         (rx_is_lockedtoref),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //   rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata        (rx_is_lockedtodata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  rx_is_lockedtodata.rx_is_lockedtodata
		.tx_std_coreclkin          (tx_std_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    tx_std_coreclkin.tx_std_coreclkin
		.rx_std_coreclkin          (rx_std_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    rx_std_coreclkin.rx_std_coreclkin
		.tx_std_clkout             (tx_std_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       tx_std_clkout.tx_std_clkout
		.rx_std_clkout             (rx_std_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       rx_std_clkout.rx_std_clkout
		.tx_std_elecidle           (tx_std_elecidle),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     tx_std_elecidle.tx_std_elecidle
		.rx_std_signaldetect       (rx_std_signaldetect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // rx_std_signaldetect.rx_std_signaldetect
		.tx_cal_busy               (tx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         rx_cal_busy.rx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  reconfig_from_xcvr.reconfig_from_xcvr
		.tx_parallel_data          ({unused_tx_parallel_data[7],unused_tx_parallel_data[6],tx_datak[3],tx_parallel_data[31],tx_parallel_data[30],tx_parallel_data[29],tx_parallel_data[28],tx_parallel_data[27],tx_parallel_data[26],tx_parallel_data[25],tx_parallel_data[24],unused_tx_parallel_data[5],unused_tx_parallel_data[4],tx_datak[2],tx_parallel_data[23],tx_parallel_data[22],tx_parallel_data[21],tx_parallel_data[20],tx_parallel_data[19],tx_parallel_data[18],tx_parallel_data[17],tx_parallel_data[16],unused_tx_parallel_data[3],unused_tx_parallel_data[2],tx_datak[1],tx_parallel_data[15],tx_parallel_data[14],tx_parallel_data[13],tx_parallel_data[12],tx_parallel_data[11],tx_parallel_data[10],tx_parallel_data[9],tx_parallel_data[8],unused_tx_parallel_data[1],unused_tx_parallel_data[0],tx_datak[0],tx_parallel_data[7],tx_parallel_data[6],tx_parallel_data[5],tx_parallel_data[4],tx_parallel_data[3],tx_parallel_data[2],tx_parallel_data[1],tx_parallel_data[0]}),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //    tx_parallel_data.tx_parallel_data
		.rx_parallel_data          ({av_sata_xcvr_core_inst_rx_parallel_data[63],av_sata_xcvr_core_inst_rx_parallel_data[62],av_sata_xcvr_core_inst_rx_parallel_data[61],av_sata_xcvr_core_inst_rx_parallel_data[60],av_sata_xcvr_core_inst_rx_parallel_data[59],av_sata_xcvr_core_inst_rx_parallel_data[58],av_sata_xcvr_core_inst_rx_parallel_data[57],av_sata_xcvr_core_inst_rx_parallel_data[56],av_sata_xcvr_core_inst_rx_parallel_data[55],av_sata_xcvr_core_inst_rx_parallel_data[54],av_sata_xcvr_core_inst_rx_parallel_data[53],av_sata_xcvr_core_inst_rx_parallel_data[52],av_sata_xcvr_core_inst_rx_parallel_data[51],av_sata_xcvr_core_inst_rx_parallel_data[50],av_sata_xcvr_core_inst_rx_parallel_data[49],av_sata_xcvr_core_inst_rx_parallel_data[48],av_sata_xcvr_core_inst_rx_parallel_data[47],av_sata_xcvr_core_inst_rx_parallel_data[46],av_sata_xcvr_core_inst_rx_parallel_data[45],av_sata_xcvr_core_inst_rx_parallel_data[44],av_sata_xcvr_core_inst_rx_parallel_data[43],av_sata_xcvr_core_inst_rx_parallel_data[42],av_sata_xcvr_core_inst_rx_parallel_data[41],av_sata_xcvr_core_inst_rx_parallel_data[40],av_sata_xcvr_core_inst_rx_parallel_data[39],av_sata_xcvr_core_inst_rx_parallel_data[38],av_sata_xcvr_core_inst_rx_parallel_data[37],av_sata_xcvr_core_inst_rx_parallel_data[36],av_sata_xcvr_core_inst_rx_parallel_data[35],av_sata_xcvr_core_inst_rx_parallel_data[34],av_sata_xcvr_core_inst_rx_parallel_data[33],av_sata_xcvr_core_inst_rx_parallel_data[32],av_sata_xcvr_core_inst_rx_parallel_data[31],av_sata_xcvr_core_inst_rx_parallel_data[30],av_sata_xcvr_core_inst_rx_parallel_data[29],av_sata_xcvr_core_inst_rx_parallel_data[28],av_sata_xcvr_core_inst_rx_parallel_data[27],av_sata_xcvr_core_inst_rx_parallel_data[26],av_sata_xcvr_core_inst_rx_parallel_data[25],av_sata_xcvr_core_inst_rx_parallel_data[24],av_sata_xcvr_core_inst_rx_parallel_data[23],av_sata_xcvr_core_inst_rx_parallel_data[22],av_sata_xcvr_core_inst_rx_parallel_data[21],av_sata_xcvr_core_inst_rx_parallel_data[20],av_sata_xcvr_core_inst_rx_parallel_data[19],av_sata_xcvr_core_inst_rx_parallel_data[18],av_sata_xcvr_core_inst_rx_parallel_data[17],av_sata_xcvr_core_inst_rx_parallel_data[16],av_sata_xcvr_core_inst_rx_parallel_data[15],av_sata_xcvr_core_inst_rx_parallel_data[14],av_sata_xcvr_core_inst_rx_parallel_data[13],av_sata_xcvr_core_inst_rx_parallel_data[12],av_sata_xcvr_core_inst_rx_parallel_data[11],av_sata_xcvr_core_inst_rx_parallel_data[10],av_sata_xcvr_core_inst_rx_parallel_data[9],av_sata_xcvr_core_inst_rx_parallel_data[8],av_sata_xcvr_core_inst_rx_parallel_data[7],av_sata_xcvr_core_inst_rx_parallel_data[6],av_sata_xcvr_core_inst_rx_parallel_data[5],av_sata_xcvr_core_inst_rx_parallel_data[4],av_sata_xcvr_core_inst_rx_parallel_data[3],av_sata_xcvr_core_inst_rx_parallel_data[2],av_sata_xcvr_core_inst_rx_parallel_data[1],av_sata_xcvr_core_inst_rx_parallel_data[0]}), //    rx_parallel_data.rx_parallel_data
		.tx_pll_refclk             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_pma_parallel_data      (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.pll_locked                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_parallel_data      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_clkslip                (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_clklow                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_fref                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_set_locktodata         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_set_locktoref          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_seriallpbken           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_signaldetect           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_prbs_done          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_prbs_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_std_pcfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_std_pcfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_pcfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_pcfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_byteorder_ena      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_byteorder_flag     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_rmfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_rmfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_wa_patternalign    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rx_std_bitslipboundarysel (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_bitslip            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_runlength_err      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_bitrev_ena         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_byterev_ena        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_std_polinv             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_polinv             (1'b0)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
	);

	assign rx_patterndetect = { av_sata_xcvr_core_inst_rx_parallel_data[60], av_sata_xcvr_core_inst_rx_parallel_data[44], av_sata_xcvr_core_inst_rx_parallel_data[28], av_sata_xcvr_core_inst_rx_parallel_data[12] };

	assign rx_runningdisp = { av_sata_xcvr_core_inst_rx_parallel_data[63], av_sata_xcvr_core_inst_rx_parallel_data[47], av_sata_xcvr_core_inst_rx_parallel_data[31], av_sata_xcvr_core_inst_rx_parallel_data[15] };

	assign rx_disperr = { av_sata_xcvr_core_inst_rx_parallel_data[59], av_sata_xcvr_core_inst_rx_parallel_data[43], av_sata_xcvr_core_inst_rx_parallel_data[27], av_sata_xcvr_core_inst_rx_parallel_data[11] };

	assign unused_rx_parallel_data = { av_sata_xcvr_core_inst_rx_parallel_data[62], av_sata_xcvr_core_inst_rx_parallel_data[61], av_sata_xcvr_core_inst_rx_parallel_data[46], av_sata_xcvr_core_inst_rx_parallel_data[45], av_sata_xcvr_core_inst_rx_parallel_data[30], av_sata_xcvr_core_inst_rx_parallel_data[29], av_sata_xcvr_core_inst_rx_parallel_data[14], av_sata_xcvr_core_inst_rx_parallel_data[13] };

	assign rx_parallel_data = { av_sata_xcvr_core_inst_rx_parallel_data[55], av_sata_xcvr_core_inst_rx_parallel_data[54], av_sata_xcvr_core_inst_rx_parallel_data[53], av_sata_xcvr_core_inst_rx_parallel_data[52], av_sata_xcvr_core_inst_rx_parallel_data[51], av_sata_xcvr_core_inst_rx_parallel_data[50], av_sata_xcvr_core_inst_rx_parallel_data[49], av_sata_xcvr_core_inst_rx_parallel_data[48], av_sata_xcvr_core_inst_rx_parallel_data[39], av_sata_xcvr_core_inst_rx_parallel_data[38], av_sata_xcvr_core_inst_rx_parallel_data[37], av_sata_xcvr_core_inst_rx_parallel_data[36], av_sata_xcvr_core_inst_rx_parallel_data[35], av_sata_xcvr_core_inst_rx_parallel_data[34], av_sata_xcvr_core_inst_rx_parallel_data[33], av_sata_xcvr_core_inst_rx_parallel_data[32], av_sata_xcvr_core_inst_rx_parallel_data[23], av_sata_xcvr_core_inst_rx_parallel_data[22], av_sata_xcvr_core_inst_rx_parallel_data[21], av_sata_xcvr_core_inst_rx_parallel_data[20], av_sata_xcvr_core_inst_rx_parallel_data[19], av_sata_xcvr_core_inst_rx_parallel_data[18], av_sata_xcvr_core_inst_rx_parallel_data[17], av_sata_xcvr_core_inst_rx_parallel_data[16], av_sata_xcvr_core_inst_rx_parallel_data[7], av_sata_xcvr_core_inst_rx_parallel_data[6], av_sata_xcvr_core_inst_rx_parallel_data[5], av_sata_xcvr_core_inst_rx_parallel_data[4], av_sata_xcvr_core_inst_rx_parallel_data[3], av_sata_xcvr_core_inst_rx_parallel_data[2], av_sata_xcvr_core_inst_rx_parallel_data[1], av_sata_xcvr_core_inst_rx_parallel_data[0] };

	assign rx_errdetect = { av_sata_xcvr_core_inst_rx_parallel_data[57], av_sata_xcvr_core_inst_rx_parallel_data[41], av_sata_xcvr_core_inst_rx_parallel_data[25], av_sata_xcvr_core_inst_rx_parallel_data[9] };

	assign rx_datak = { av_sata_xcvr_core_inst_rx_parallel_data[56], av_sata_xcvr_core_inst_rx_parallel_data[40], av_sata_xcvr_core_inst_rx_parallel_data[24], av_sata_xcvr_core_inst_rx_parallel_data[8] };

	assign rx_syncstatus = { av_sata_xcvr_core_inst_rx_parallel_data[58], av_sata_xcvr_core_inst_rx_parallel_data[42], av_sata_xcvr_core_inst_rx_parallel_data[26], av_sata_xcvr_core_inst_rx_parallel_data[10] };

endmodule
