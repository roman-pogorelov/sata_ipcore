// megafunction wizard: %Stratix V Transceiver Native PHY v17.1%
// GENERATION: XML
// sv_sata_xcvr_core.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module sv_sata_xcvr_core (
		input  wire [0:0]  pll_powerdown,           //           pll_powerdown.pll_powerdown
		input  wire [0:0]  tx_analogreset,          //          tx_analogreset.tx_analogreset
		input  wire [0:0]  tx_digitalreset,         //         tx_digitalreset.tx_digitalreset
		output wire [0:0]  tx_serial_data,          //          tx_serial_data.tx_serial_data
		input  wire [0:0]  ext_pll_clk,             //             ext_pll_clk.ext_pll_clk
		input  wire [0:0]  rx_analogreset,          //          rx_analogreset.rx_analogreset
		input  wire [0:0]  rx_digitalreset,         //         rx_digitalreset.rx_digitalreset
		input  wire [0:0]  rx_cdr_refclk,           //           rx_cdr_refclk.rx_cdr_refclk
		input  wire [0:0]  rx_serial_data,          //          rx_serial_data.rx_serial_data
		output wire [0:0]  rx_is_lockedtoref,       //       rx_is_lockedtoref.rx_is_lockedtoref
		output wire [0:0]  rx_is_lockedtodata,      //      rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [0:0]  tx_std_coreclkin,        //        tx_std_coreclkin.tx_std_coreclkin
		input  wire [0:0]  rx_std_coreclkin,        //        rx_std_coreclkin.rx_std_coreclkin
		output wire [0:0]  tx_std_clkout,           //           tx_std_clkout.tx_std_clkout
		output wire [0:0]  rx_std_clkout,           //           rx_std_clkout.rx_std_clkout
		input  wire [0:0]  tx_std_elecidle,         //         tx_std_elecidle.tx_std_elecidle
		output wire [0:0]  rx_std_signaldetect,     //     rx_std_signaldetect.rx_std_signaldetect
		output wire [0:0]  tx_cal_busy,             //             tx_cal_busy.tx_cal_busy
		output wire [0:0]  rx_cal_busy,             //             rx_cal_busy.rx_cal_busy
		input  wire [69:0] reconfig_to_xcvr,        //        reconfig_to_xcvr.reconfig_to_xcvr
		output wire [45:0] reconfig_from_xcvr,      //      reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [31:0] tx_parallel_data,        //        tx_parallel_data.tx_parallel_data
		input  wire [3:0]  tx_datak,                //                tx_datak.tx_datak
		input  wire [27:0] unused_tx_parallel_data, // unused_tx_parallel_data.unused_tx_parallel_data
		output wire [31:0] rx_parallel_data,        //        rx_parallel_data.rx_parallel_data
		output wire [3:0]  rx_datak,                //                rx_datak.rx_datak
		output wire [3:0]  rx_errdetect,            //            rx_errdetect.rx_errdetect
		output wire [3:0]  rx_disperr,              //              rx_disperr.rx_disperr
		output wire [3:0]  rx_runningdisp,          //          rx_runningdisp.rx_runningdisp
		output wire [3:0]  rx_patterndetect,        //        rx_patterndetect.rx_patterndetect
		output wire [3:0]  rx_syncstatus,           //           rx_syncstatus.rx_syncstatus
		output wire [7:0]  unused_rx_parallel_data  // unused_rx_parallel_data.unused_rx_parallel_data
	);

	wire  [63:0] sv_sata_xcvr_core_inst_rx_parallel_data; // port fragment

	altera_xcvr_native_sv #(
		.tx_enable                       (1),
		.rx_enable                       (1),
		.enable_std                      (1),
		.enable_teng                     (0),
		.data_path_select                ("standard"),
		.channels                        (1),
		.bonded_mode                     ("non_bonded"),
		.data_rate                       ("6000 Mbps"),
		.pma_width                       (20),
		.tx_pma_clk_div                  (1),
		.tx_pma_txdetectrx_ctrl          (0),
		.pll_reconfig_enable             (0),
		.pll_external_enable             (1),
		.pll_data_rate                   ("6000 Mbps"),
		.pll_type                        ("CMU"),
		.pll_network_select              ("x1"),
		.plls                            (1),
		.pll_select                      (0),
		.pll_refclk_cnt                  (1),
		.pll_refclk_select               ("0"),
		.pll_refclk_freq                 ("125.0 MHz"),
		.pll_feedback_path               ("internal"),
		.cdr_reconfig_enable             (0),
		.cdr_refclk_cnt                  (1),
		.cdr_refclk_select               (0),
		.cdr_refclk_freq                 ("150.0 MHz"),
		.rx_ppm_detect_threshold         ("1000"),
		.rx_clkslip_enable               (0),
		.std_protocol_hint               ("basic"),
		.std_pcs_pma_width               (20),
		.std_low_latency_bypass_enable   (0),
		.std_tx_pcfifo_mode              ("low_latency"),
		.std_rx_pcfifo_mode              ("low_latency"),
		.std_rx_byte_order_enable        (0),
		.std_rx_byte_order_mode          ("manual"),
		.std_rx_byte_order_width         (9),
		.std_rx_byte_order_symbol_count  (1),
		.std_rx_byte_order_pattern       ("0"),
		.std_rx_byte_order_pad           ("0"),
		.std_tx_byte_ser_enable          (1),
		.std_rx_byte_deser_enable        (1),
		.std_tx_8b10b_enable             (1),
		.std_tx_8b10b_disp_ctrl_enable   (0),
		.std_rx_8b10b_enable             (1),
		.std_rx_rmfifo_enable            (0),
		.std_rx_rmfifo_pattern_p         ("00000"),
		.std_rx_rmfifo_pattern_n         ("00000"),
		.std_tx_bitslip_enable           (0),
		.std_rx_word_aligner_mode        ("manual"),
		.std_rx_word_aligner_pattern_len (10),
		.std_rx_word_aligner_pattern     ("17c"),
		.std_rx_word_aligner_rknumber    (3),
		.std_rx_word_aligner_renumber    (3),
		.std_rx_word_aligner_rgnumber    (3),
		.std_rx_run_length_val           (31),
		.std_tx_bitrev_enable            (0),
		.std_rx_bitrev_enable            (0),
		.std_tx_byterev_enable           (0),
		.std_rx_byterev_enable           (0),
		.std_tx_polinv_enable            (0),
		.std_rx_polinv_enable            (0),
		.teng_protocol_hint              ("basic"),
		.teng_pcs_pma_width              (40),
		.teng_pld_pcs_width              (40),
		.teng_txfifo_mode                ("phase_comp"),
		.teng_txfifo_full                (31),
		.teng_txfifo_empty               (0),
		.teng_txfifo_pfull               (23),
		.teng_txfifo_pempty              (2),
		.teng_rxfifo_mode                ("phase_comp"),
		.teng_rxfifo_full                (31),
		.teng_rxfifo_empty               (0),
		.teng_rxfifo_pfull               (23),
		.teng_rxfifo_pempty              (2),
		.teng_rxfifo_align_del           (0),
		.teng_rxfifo_control_del         (0),
		.teng_tx_frmgen_enable           (0),
		.teng_tx_frmgen_user_length      (2048),
		.teng_tx_frmgen_burst_enable     (0),
		.teng_rx_frmsync_enable          (0),
		.teng_rx_frmsync_user_length     (2048),
		.teng_frmgensync_diag_word       ("6400000000000000"),
		.teng_frmgensync_scrm_word       ("2800000000000000"),
		.teng_frmgensync_skip_word       ("1e1e1e1e1e1e1e1e"),
		.teng_frmgensync_sync_word       ("78f678f678f678f6"),
		.teng_tx_sh_err                  (0),
		.teng_tx_crcgen_enable           (0),
		.teng_rx_crcchk_enable           (0),
		.teng_tx_64b66b_enable           (0),
		.teng_rx_64b66b_enable           (0),
		.teng_tx_scram_enable            (0),
		.teng_tx_scram_user_seed         ("000000000000000"),
		.teng_rx_descram_enable          (0),
		.teng_tx_dispgen_enable          (0),
		.teng_rx_dispchk_enable          (0),
		.teng_rx_blksync_enable          (0),
		.teng_tx_polinv_enable           (0),
		.teng_tx_bitslip_enable          (0),
		.teng_rx_polinv_enable           (0),
		.teng_rx_bitslip_enable          (0)
	) sv_sata_xcvr_core_inst (
		.pll_powerdown             (pll_powerdown),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       pll_powerdown.pll_powerdown
		.tx_analogreset            (tx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     tx_digitalreset.tx_digitalreset
		.tx_serial_data            (tx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      tx_serial_data.tx_serial_data
		.ext_pll_clk               (ext_pll_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         ext_pll_clk.ext_pll_clk
		.rx_analogreset            (rx_analogreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      rx_analogreset.rx_analogreset
		.rx_digitalreset           (rx_digitalreset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     rx_digitalreset.rx_digitalreset
		.rx_cdr_refclk             (rx_cdr_refclk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       rx_cdr_refclk.rx_cdr_refclk
		.rx_serial_data            (rx_serial_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //      rx_serial_data.rx_serial_data
		.rx_is_lockedtoref         (rx_is_lockedtoref),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //   rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata        (rx_is_lockedtodata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  rx_is_lockedtodata.rx_is_lockedtodata
		.tx_std_coreclkin          (tx_std_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    tx_std_coreclkin.tx_std_coreclkin
		.rx_std_coreclkin          (rx_std_coreclkin),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    rx_std_coreclkin.rx_std_coreclkin
		.tx_std_clkout             (tx_std_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       tx_std_clkout.tx_std_clkout
		.rx_std_clkout             (rx_std_clkout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       rx_std_clkout.rx_std_clkout
		.tx_std_elecidle           (tx_std_elecidle),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     tx_std_elecidle.tx_std_elecidle
		.rx_std_signaldetect       (rx_std_signaldetect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // rx_std_signaldetect.rx_std_signaldetect
		.tx_cal_busy               (tx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         rx_cal_busy.rx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //  reconfig_from_xcvr.reconfig_from_xcvr
		.tx_parallel_data          ({unused_tx_parallel_data[27],unused_tx_parallel_data[26],unused_tx_parallel_data[25],unused_tx_parallel_data[24],unused_tx_parallel_data[23],unused_tx_parallel_data[22],unused_tx_parallel_data[21],unused_tx_parallel_data[20],unused_tx_parallel_data[19],unused_tx_parallel_data[18],unused_tx_parallel_data[17],unused_tx_parallel_data[16],unused_tx_parallel_data[15],unused_tx_parallel_data[14],unused_tx_parallel_data[13],unused_tx_parallel_data[12],unused_tx_parallel_data[11],unused_tx_parallel_data[10],unused_tx_parallel_data[9],unused_tx_parallel_data[8],unused_tx_parallel_data[7],unused_tx_parallel_data[6],tx_datak[3],tx_parallel_data[31],tx_parallel_data[30],tx_parallel_data[29],tx_parallel_data[28],tx_parallel_data[27],tx_parallel_data[26],tx_parallel_data[25],tx_parallel_data[24],unused_tx_parallel_data[5],unused_tx_parallel_data[4],tx_datak[2],tx_parallel_data[23],tx_parallel_data[22],tx_parallel_data[21],tx_parallel_data[20],tx_parallel_data[19],tx_parallel_data[18],tx_parallel_data[17],tx_parallel_data[16],unused_tx_parallel_data[3],unused_tx_parallel_data[2],tx_datak[1],tx_parallel_data[15],tx_parallel_data[14],tx_parallel_data[13],tx_parallel_data[12],tx_parallel_data[11],tx_parallel_data[10],tx_parallel_data[9],tx_parallel_data[8],unused_tx_parallel_data[1],unused_tx_parallel_data[0],tx_datak[0],tx_parallel_data[7],tx_parallel_data[6],tx_parallel_data[5],tx_parallel_data[4],tx_parallel_data[3],tx_parallel_data[2],tx_parallel_data[1],tx_parallel_data[0]}),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //    tx_parallel_data.tx_parallel_data
		.rx_parallel_data          ({sv_sata_xcvr_core_inst_rx_parallel_data[63],sv_sata_xcvr_core_inst_rx_parallel_data[62],sv_sata_xcvr_core_inst_rx_parallel_data[61],sv_sata_xcvr_core_inst_rx_parallel_data[60],sv_sata_xcvr_core_inst_rx_parallel_data[59],sv_sata_xcvr_core_inst_rx_parallel_data[58],sv_sata_xcvr_core_inst_rx_parallel_data[57],sv_sata_xcvr_core_inst_rx_parallel_data[56],sv_sata_xcvr_core_inst_rx_parallel_data[55],sv_sata_xcvr_core_inst_rx_parallel_data[54],sv_sata_xcvr_core_inst_rx_parallel_data[53],sv_sata_xcvr_core_inst_rx_parallel_data[52],sv_sata_xcvr_core_inst_rx_parallel_data[51],sv_sata_xcvr_core_inst_rx_parallel_data[50],sv_sata_xcvr_core_inst_rx_parallel_data[49],sv_sata_xcvr_core_inst_rx_parallel_data[48],sv_sata_xcvr_core_inst_rx_parallel_data[47],sv_sata_xcvr_core_inst_rx_parallel_data[46],sv_sata_xcvr_core_inst_rx_parallel_data[45],sv_sata_xcvr_core_inst_rx_parallel_data[44],sv_sata_xcvr_core_inst_rx_parallel_data[43],sv_sata_xcvr_core_inst_rx_parallel_data[42],sv_sata_xcvr_core_inst_rx_parallel_data[41],sv_sata_xcvr_core_inst_rx_parallel_data[40],sv_sata_xcvr_core_inst_rx_parallel_data[39],sv_sata_xcvr_core_inst_rx_parallel_data[38],sv_sata_xcvr_core_inst_rx_parallel_data[37],sv_sata_xcvr_core_inst_rx_parallel_data[36],sv_sata_xcvr_core_inst_rx_parallel_data[35],sv_sata_xcvr_core_inst_rx_parallel_data[34],sv_sata_xcvr_core_inst_rx_parallel_data[33],sv_sata_xcvr_core_inst_rx_parallel_data[32],sv_sata_xcvr_core_inst_rx_parallel_data[31],sv_sata_xcvr_core_inst_rx_parallel_data[30],sv_sata_xcvr_core_inst_rx_parallel_data[29],sv_sata_xcvr_core_inst_rx_parallel_data[28],sv_sata_xcvr_core_inst_rx_parallel_data[27],sv_sata_xcvr_core_inst_rx_parallel_data[26],sv_sata_xcvr_core_inst_rx_parallel_data[25],sv_sata_xcvr_core_inst_rx_parallel_data[24],sv_sata_xcvr_core_inst_rx_parallel_data[23],sv_sata_xcvr_core_inst_rx_parallel_data[22],sv_sata_xcvr_core_inst_rx_parallel_data[21],sv_sata_xcvr_core_inst_rx_parallel_data[20],sv_sata_xcvr_core_inst_rx_parallel_data[19],sv_sata_xcvr_core_inst_rx_parallel_data[18],sv_sata_xcvr_core_inst_rx_parallel_data[17],sv_sata_xcvr_core_inst_rx_parallel_data[16],sv_sata_xcvr_core_inst_rx_parallel_data[15],sv_sata_xcvr_core_inst_rx_parallel_data[14],sv_sata_xcvr_core_inst_rx_parallel_data[13],sv_sata_xcvr_core_inst_rx_parallel_data[12],sv_sata_xcvr_core_inst_rx_parallel_data[11],sv_sata_xcvr_core_inst_rx_parallel_data[10],sv_sata_xcvr_core_inst_rx_parallel_data[9],sv_sata_xcvr_core_inst_rx_parallel_data[8],sv_sata_xcvr_core_inst_rx_parallel_data[7],sv_sata_xcvr_core_inst_rx_parallel_data[6],sv_sata_xcvr_core_inst_rx_parallel_data[5],sv_sata_xcvr_core_inst_rx_parallel_data[4],sv_sata_xcvr_core_inst_rx_parallel_data[3],sv_sata_xcvr_core_inst_rx_parallel_data[2],sv_sata_xcvr_core_inst_rx_parallel_data[1],sv_sata_xcvr_core_inst_rx_parallel_data[0]}), //    rx_parallel_data.rx_parallel_data
		.tx_pll_refclk             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_pma_pclk               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_pma_parallel_data      (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.pll_locked                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_pclk               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_parallel_data      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_clkslip                (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_clklow                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_fref                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_set_locktodata         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_set_locktoref          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_seriallpbken           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_signaldetect           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_pma_qpipulldn          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_qpipullup          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_qpipulldn          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_txdetectrx         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_pma_rxfound            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_prbs_done          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_prbs_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_std_pcfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_std_pcfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_pcfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_pcfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_byteorder_ena      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_byteorder_flag     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_rmfifo_full        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_rmfifo_empty       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_wa_patternalign    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rx_std_bitslipboundarysel (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_bitslip            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_runlength_err      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_std_bitrev_ena         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_byterev_ena        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_std_polinv             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_std_polinv             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_10g_coreclkin          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_coreclkin          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_10g_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_clkout             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_clk33out           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_prbs_err_clr       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_prbs_done          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_prbs_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_control            (9'b000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rx_10g_control            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_data_valid         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_10g_fifo_full          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_fifo_pfull         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_fifo_empty         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_fifo_pempty        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_fifo_del           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_fifo_insert        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_rd_en         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_data_valid         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_full          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_pfull         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_empty         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_pempty        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_del           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_insert        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_align_val     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_fifo_align_clr     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_fifo_align_en      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.tx_10g_frame              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_frame_diag_status  (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //         (terminated)
		.tx_10g_frame_burst_en     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_frame              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_lock         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_mfrm_err     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_sync_err     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_skip_ins     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_pyld_ins     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_skip_err     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_diag_err     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_frame_diag_status  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_crc32_err          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_descram_err        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_blk_lock           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_blk_sh_err         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.tx_10g_bitslip            (7'b0000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //         (terminated)
		.rx_10g_bitslip            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_highber            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //         (terminated)
		.rx_10g_highber_clr_cnt    (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         (terminated)
		.rx_10g_clr_errblk_count   (1'b0)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
	);

	assign rx_parallel_data = { sv_sata_xcvr_core_inst_rx_parallel_data[55], sv_sata_xcvr_core_inst_rx_parallel_data[54], sv_sata_xcvr_core_inst_rx_parallel_data[53], sv_sata_xcvr_core_inst_rx_parallel_data[52], sv_sata_xcvr_core_inst_rx_parallel_data[51], sv_sata_xcvr_core_inst_rx_parallel_data[50], sv_sata_xcvr_core_inst_rx_parallel_data[49], sv_sata_xcvr_core_inst_rx_parallel_data[48], sv_sata_xcvr_core_inst_rx_parallel_data[39], sv_sata_xcvr_core_inst_rx_parallel_data[38], sv_sata_xcvr_core_inst_rx_parallel_data[37], sv_sata_xcvr_core_inst_rx_parallel_data[36], sv_sata_xcvr_core_inst_rx_parallel_data[35], sv_sata_xcvr_core_inst_rx_parallel_data[34], sv_sata_xcvr_core_inst_rx_parallel_data[33], sv_sata_xcvr_core_inst_rx_parallel_data[32], sv_sata_xcvr_core_inst_rx_parallel_data[23], sv_sata_xcvr_core_inst_rx_parallel_data[22], sv_sata_xcvr_core_inst_rx_parallel_data[21], sv_sata_xcvr_core_inst_rx_parallel_data[20], sv_sata_xcvr_core_inst_rx_parallel_data[19], sv_sata_xcvr_core_inst_rx_parallel_data[18], sv_sata_xcvr_core_inst_rx_parallel_data[17], sv_sata_xcvr_core_inst_rx_parallel_data[16], sv_sata_xcvr_core_inst_rx_parallel_data[7], sv_sata_xcvr_core_inst_rx_parallel_data[6], sv_sata_xcvr_core_inst_rx_parallel_data[5], sv_sata_xcvr_core_inst_rx_parallel_data[4], sv_sata_xcvr_core_inst_rx_parallel_data[3], sv_sata_xcvr_core_inst_rx_parallel_data[2], sv_sata_xcvr_core_inst_rx_parallel_data[1], sv_sata_xcvr_core_inst_rx_parallel_data[0] };

	assign rx_disperr = { sv_sata_xcvr_core_inst_rx_parallel_data[59], sv_sata_xcvr_core_inst_rx_parallel_data[43], sv_sata_xcvr_core_inst_rx_parallel_data[27], sv_sata_xcvr_core_inst_rx_parallel_data[11] };

	assign rx_runningdisp = { sv_sata_xcvr_core_inst_rx_parallel_data[63], sv_sata_xcvr_core_inst_rx_parallel_data[47], sv_sata_xcvr_core_inst_rx_parallel_data[31], sv_sata_xcvr_core_inst_rx_parallel_data[15] };

	assign rx_patterndetect = { sv_sata_xcvr_core_inst_rx_parallel_data[60], sv_sata_xcvr_core_inst_rx_parallel_data[44], sv_sata_xcvr_core_inst_rx_parallel_data[28], sv_sata_xcvr_core_inst_rx_parallel_data[12] };

	assign rx_syncstatus = { sv_sata_xcvr_core_inst_rx_parallel_data[58], sv_sata_xcvr_core_inst_rx_parallel_data[42], sv_sata_xcvr_core_inst_rx_parallel_data[26], sv_sata_xcvr_core_inst_rx_parallel_data[10] };

	assign rx_errdetect = { sv_sata_xcvr_core_inst_rx_parallel_data[57], sv_sata_xcvr_core_inst_rx_parallel_data[41], sv_sata_xcvr_core_inst_rx_parallel_data[25], sv_sata_xcvr_core_inst_rx_parallel_data[9] };

	assign unused_rx_parallel_data = { sv_sata_xcvr_core_inst_rx_parallel_data[62], sv_sata_xcvr_core_inst_rx_parallel_data[61], sv_sata_xcvr_core_inst_rx_parallel_data[46], sv_sata_xcvr_core_inst_rx_parallel_data[45], sv_sata_xcvr_core_inst_rx_parallel_data[30], sv_sata_xcvr_core_inst_rx_parallel_data[29], sv_sata_xcvr_core_inst_rx_parallel_data[14], sv_sata_xcvr_core_inst_rx_parallel_data[13] };

	assign rx_datak = { sv_sata_xcvr_core_inst_rx_parallel_data[56], sv_sata_xcvr_core_inst_rx_parallel_data[40], sv_sata_xcvr_core_inst_rx_parallel_data[24], sv_sata_xcvr_core_inst_rx_parallel_data[8] };

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_native_sv" version="17.1" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="show_advanced_features" value="0" />
// Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
// Retrieval info: 	<generic name="message_level" value="error" />
// Retrieval info: 	<generic name="tx_enable" value="1" />
// Retrieval info: 	<generic name="rx_enable" value="1" />
// Retrieval info: 	<generic name="enable_std" value="1" />
// Retrieval info: 	<generic name="enable_teng" value="0" />
// Retrieval info: 	<generic name="set_data_path_select" value="standard" />
// Retrieval info: 	<generic name="channels" value="1" />
// Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
// Retrieval info: 	<generic name="enable_simple_interface" value="1" />
// Retrieval info: 	<generic name="set_data_rate" value="6000" />
// Retrieval info: 	<generic name="pma_direct_width" value="80" />
// Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
// Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
// Retrieval info: 	<generic name="pll_external_enable" value="1" />
// Retrieval info: 	<generic name="plls" value="1" />
// Retrieval info: 	<generic name="pll_select" value="0" />
// Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
// Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
// Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
// Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
// Retrieval info: 	<generic name="set_cdr_refclk_freq" value="150.0 MHz" />
// Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
// Retrieval info: 	<generic name="enable_port_tx_pma_qpipullup" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_qpipulldn" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_txdetectrx" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_rxfound" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_pclk" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_pma_qpipulldn" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_pma_pclk" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
// Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
// Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="0" />
// Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
// Retrieval info: 	<generic name="std_pcs_pma_width" value="20" />
// Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
// Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="low_latency" />
// Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
// Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
// Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
// Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
// Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
// Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="1" />
// Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="1" />
// Retrieval info: 	<generic name="std_tx_8b10b_enable" value="1" />
// Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_8b10b_enable" value="1" />
// Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
// Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
// Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
// Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
// Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="manual" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="10" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="17c" />
// Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
// Retrieval info: 	<generic name="std_rx_run_length_val" value="31" />
// Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
// Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
// Retrieval info: 	<generic name="teng_protocol_hint" value="basic" />
// Retrieval info: 	<generic name="teng_pcs_pma_width" value="40" />
// Retrieval info: 	<generic name="teng_pld_pcs_width" value="40" />
// Retrieval info: 	<generic name="teng_txfifo_mode" value="phase_comp" />
// Retrieval info: 	<generic name="teng_txfifo_full" value="31" />
// Retrieval info: 	<generic name="teng_txfifo_empty" value="0" />
// Retrieval info: 	<generic name="teng_txfifo_pfull" value="23" />
// Retrieval info: 	<generic name="teng_txfifo_pempty" value="2" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pfull" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_empty" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pempty" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_del" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_fifo_insert" value="0" />
// Retrieval info: 	<generic name="teng_rxfifo_mode" value="phase_comp" />
// Retrieval info: 	<generic name="teng_rxfifo_full" value="31" />
// Retrieval info: 	<generic name="teng_rxfifo_empty" value="0" />
// Retrieval info: 	<generic name="teng_rxfifo_pfull" value="23" />
// Retrieval info: 	<generic name="teng_rxfifo_pempty" value="2" />
// Retrieval info: 	<generic name="teng_rxfifo_align_del" value="0" />
// Retrieval info: 	<generic name="teng_rxfifo_control_del" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_data_valid" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pfull" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_empty" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pempty" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_del" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_insert" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_rd_en" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_val" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_clr" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_en" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_clk33out" value="0" />
// Retrieval info: 	<generic name="teng_tx_frmgen_user_length" value="2048" />
// Retrieval info: 	<generic name="teng_tx_frmgen_burst_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_frame" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_frame_diag_status" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_frame_burst_en" value="0" />
// Retrieval info: 	<generic name="teng_rx_frmsync_user_length" value="2048" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_lock" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_mfrm_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_sync_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_pyld_ins" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_ins" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_status" value="0" />
// Retrieval info: 	<generic name="teng_tx_sh_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_crc32_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_highber" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_highber_clr_cnt" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_clr_errblk_count" value="0" />
// Retrieval info: 	<generic name="teng_tx_scram_user_seed" value="000000000000000" />
// Retrieval info: 	<generic name="enable_port_rx_10g_descram_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_blk_lock" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_blk_sh_err" value="0" />
// Retrieval info: 	<generic name="teng_tx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="teng_tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="teng_rx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="teng_rx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_10g_bitslip" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_10g_bitslip" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_teng_prbs_status" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : sv_sata_xcvr_core.vo
// RELATED_FILES: sv_sata_xcvr_core.v, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_native_sv_functions_h.sv, altera_xcvr_native_sv.sv
