// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:01:49 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P+JHLbOPel0YaeFd2xZsuMhU5cM/nOfjeNo9dRIVmZlPl8QHrmRwM2howwQNd/yJ
aJpdMlcEp6gu6EGGdvmka/yBVPo7WuAGtlMYjOztOsscNurkycE2swmAuT4usQAZ
KNVy5DMZ3fV83TqRHd72ErUS1YyFO/QG+QXVYnsiycg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48656)
k0lwjQyT7u8PFVxTHqyLQpwyL1pFi7KNkDWWcqbBB++jML5H8M5m986n6gRI5FJb
A0z8FOXbCYSU5RJmuDrME+mTX/uQrqFn7N8OsD1O2tZiLSdS8yqh0b9WZl4Xmrz3
AskMWI7EyeGcK7raCy5P4Q38p4UulqDTPVSATzSwhRbiR/Nd2ikiPII7IRGuscED
kMEKsLhDi6l5wPyZw6bDpKAYTCgFTclUJ4fNGGCck/4GBJIU3pSBgwRH8u467kYi
Qp4HwWgKL0kc9q7bFYs1IkWTnfxhbME8HGqks9PXhdQXm9G6/ieES5bcwYBRd8Kp
nDvmVyvqGpOlEYmUgzRciHkliE1Q43A1Og1LNRF4obCPtYyQ0ZE+yMPDCEyPc/HF
SL2vqiAaxY343AfqGJTIfjV5DgeUNlYq6jZpFqE1YrBR1uCw9TKP1ARkymLf0Gi/
yGas8QvfrHvjIn+YSk0+r0KzbTlr6LKiS8H8YeiMx3Fy8kWHErSMJMPSpqPOUCyr
fuwBdE71hS4UNwQiqICkj7k62PdddAg/XtkP7QqsUSTG7f1ldmw/q4s0egT3ImtB
HtAdqyGOxsueGIv+Pbj0ORbTiXNVd1hJRWkJ8x8rB4A1OKFUKLdjAJqZ6jX7AcVu
/xzl4zopAi+WWY1dDxXTcd/6pRgm8Zi01H6nD93oaABKCFnR1Qr+v/D3nYMlk1vl
tmmoh+jlJZQTsHjc2NxAd+ZN1j33BLknVVwWBiGF6SQ+cZHs6Hj7L1CQJ9iRMM/N
8Ze85yKAAXb8akBkHD9FhYeKl0PfPK+ksFW3BhqJa8dRa2iKktDdJ7P861jo1EA1
k2Z55y+QcKzd07Pi/1x3ubfhewtuJTolrQQtWUz2+rGz4hW0sE/SWYJEyFnuuphu
RNZrefFib/4sRf7a99AwjSy8zlJWvQ3T/cbf16kOUOiWiB4+/NAlrKXx2/UviMyM
wjYnI/rrhKgy+YkH0LqRbDLC4SACGUakxeo3wuBT6mBBLRzNUoT1h+yMX6r/U7Zb
o3SA0sQXY1iPiXEOXqLKRSIgNRU39MXcxwkQH2N+xTsUYWolllVrtqcX/EutZqsd
M3L9n2xILrUeyRpJqwyvW3O1bt7QiIyhjyukk1HLq/9JGVoNkPI9GlawgnceJUcI
j58uME+YdNJTMVJgXh1FBYP5XiSdDb6jdXB8NGBC7k/zgAkB9pP+bMrDOr4GeA7x
06kPVEm2CGpY/B7f6JxD9egcReBLGOgbQ8k/ObK8WQ2xhu6t0tN+6Nu9AvWJQoUI
4SzhwDDtkyxUcQO3On9mjTVKQhIo0xzmQ2JUJ1jPJpM2MQ7TmnFiGhJ8t9ALWiA2
DAvXg+f1ffz12VuYng14yYOSRjBf07Pb3k49waZ/0TF6ICIZsPjeOe8O4S5/gWwh
YSMdrnyC3SbTT+u7mayD0EPMqQlqcUOXCOntb6dHxPkiyrpI9FvnCCQS4Zr3m5ZS
IoqWTpBQcNfCCVLOvSSM224hKB2isDbg0/2UbMQ+mvbigjb6yE/adR5P77hGERl5
7QAMAPcPKcw69GLs9+4EL95f+41Vnh5mofQbWSNj9ynWPv6WnfgBv4hPmvbhAHUx
Oji1cgGwnog/P/B4wxHeRJxuOyAyjGjbX92H2oYRfuVrkDBiCOwNhbnNh5YZDGkj
QEqN9Tu/8Nx0a3cZfKOX9SRbY1SOmA1VBmHHs9IQDizjr90hsD5EKIEPHKi9p/BY
rE46jzibJr5ai3Mgg9UCgHu/IwgH80nYPs8RKitVWFEWlDU7hT4YYE63KlWv6bgl
jN2gUUa5WwVd1+7NeAdPQOMVOlbbHfXZqMSno1yuI3L9JclzAmwuRaVZufwU63Lp
Zup0aYJEu/Qxs/wLfa5JpkpjxWxtaaUkTNkLt9b3mKNSiSTf9Ymdu1O7Cmz7aIgB
9fKwuvCAZv/nJae2IfrnOxYvZsOlGM2xB3KzJSG4f9ClumFebyn+Ls4/GNN06rL+
OukfwnnK3xLTKJtqPUn9+f5cy0KXfsUafujuZw4wlNqQpunBmYA7Hl4dKHIrXsRS
GuQIfCHMOOCxRLryULMmfJP2R60uvFbqDSO44dtmMFp1F9bz7F8ZCJHyjSQXAJUq
oE+Y2WqqH00VsVTOjRhHW4PYx/zB9X4vB7HLAJMXjXsYaIdvmjwCUXI9H/Agnxjl
4i9BjgO+Ra7ILyHMafZG7fJvpXx3dPKaSvj0hAsWuvIHirzSOL4w4F5a+P92uGXD
VCOIAoX6uxzBuMWTK7SL+6VLtDhXLL8dKtoga+Gp0a6HCDgnQSfXq1vQKnjFcOWG
HH9uKXDWBKxRAV337sZ1xifw8hHNyQD8aLrIAsJ0AnlMjGloJ6hARnm7Nq1B8OiS
xopQw0/qxMC+WlNtJ2l7AO+cuafBDc3jVKKcgEnHhvId8s3vsYqGf913QeqMzag7
fbqbv6O2tZXDMdhGpYt1Ob3+RmTw/K03kU1+X5m+9X5+DOMqK3PeKlfbK0RT4q+1
mBhj7V/9845B0TUEuxzthozrjr0P/u3dAat+T5GMZmrGwmp59kaMd9ZP+ozgQwpN
+YlWCBK6RlFxVp68ookO+cDrmoBbnhLuj39nMNr4Dm9pbLuawVHiWybwyf/KS0Oi
Y0OYjItLkM38siGnF2MsCbkxQQogPxsxAfEPoWUYR1X0DedzquaEMZJ3GMAv4r5w
NQkrA2Apk5PG4X05kGTbstZ872inlTgzjk5m7fJhQZncp42x0zAJsKWyUyZeoeyO
NvJghl9y+JYMYLu0GBNo1EKE/SITIC2HGjV7e2MZEOE+0AeIp7MUSP7Ov2B9tJ0L
UqBaLATHS4xie8RLBWrxqXeS18HAggzvn55l7gjME6Q17QyyjV7MILmHttwKwCIg
Zeg+boNP+G0Bjo7+yg1HgyRqDCyfIZG+b8NQjCVpGLOFt2QoCri7BDuL8j+xvuMV
3q3rGby3bwXQnkEYkcDCgRAyH84AhLaeSYbrE/9G4aXH1HDbvUgyLJxjphM9SNQu
9eaM8XCqmegJCcvBygeMO3CjJ7yjTE+MloP/BNCpjdh3rKIIo6DI/dEyazm70Int
6NEhzbXoQYo0T5Bx/PWQgfpD1Uu9OLdjh7naf59R3ZjYgVenWp12j0mX5uWo1sjr
l/Y18et9Tp08UvZpmAopDZfj0VNcll6eX1R7U6aAFkRmU7Z31hVg9BFZ0umMsMiA
RQwJVXG9pbgyrAn3rrTiIvT+yFTyaz9ilwf3rSIWbfBTirAGhBQMxP4UjWGacm87
K3UFbEzhPUnBrp9u75ySYls2r6xLsRSfMUA9MpZJng40UazppVyHhok0IxXnMSme
QYbO2/1/PqKmyg2TjEwJXOa9d3F5LOmWD2krx76et8s/9NR7DMM2legWiPyyln9O
jdDbeNdjXGpr3DzMVsROyLqi4Jnqhx8p6hpTQPznuxX23pY2rTiJIne8LZOXIVpe
ZLBoUoAuxIbCYyhJkEJaVzcmobTXcKAr2xCeMaW+RAerqsJl+/MaGhZQB2LMPQnj
Fs+0lw1D55GpzZulFoMdfQdoGwwEyt5eSxDRoowdDZCdukXMRhxg1MuC6h/048pK
4eoxqFhN9w1c8WGQztHLF5kcCB6Nho3+IAc7u6WUgYC/MMzdA+sa2lCAnrWxo/fH
k8qDtJMk1y1MIVcd5Q6DsTlr3Hb8tOsc8f4eYWZTTEjuNu/ofc6Hns02rjchBfPP
Z/ZfCIwQHFL2M9V5dfrB0v9OEeHh9zYv7W5GJQKB8Sfs1VXFlQsQVRx/dy2khGcQ
zuvuQLJdQnCfotEzkEgxKexiqFCybPGy/5t8Z8VRucCriEpyck9HSeBa29yhMJ9d
geqNODCFePVotB5F9Gb3F9VVs6R6E2VWl2JMAaVIfbbWz7elDfyW211mqwadL1AU
5ohC4TCBzdxV7KW1wrNJS7PRdpF8DNmJ0n3N/2tC3Py8/B+WPpEb1RyfQextxWgH
DdTQvpkU8r+V8U68BMh+nc9FtBMPdbaMIF7faxmH+yI+GM4D3to05uDpuVl5KarP
vf/7LTCbTSn4J1D6y0oSlIAfe4NFi0f50E0XI4FxDSiMhUumEIsKTzHGrCIrFGUd
LDoQGC46R9IFRDs8AKMoKfxEiGSbYfGKbk7zbvszPUtUCxjQ52eiu8W+EtjIzG9H
AMOAV4kxotWePNv8BrwLgsaUXUgtEHl/FpcqUV6obYfuwHCiE6VKPoa2cXlF5rPz
RC1se9RdsProO1fEDjnhxmtOfsEAmwjQrzMACXhO1CYk18PNUuvzMTftoUG3yaUp
mz92Y/T9J+5/gWSSsXDydVlTCjnvNq9C/l5KwsVAdiDi9ngwcUlZED+7XLddtAVV
u6RHhlnFKiaO9vzb2n4Ug33HA4jfIQpzwsPQGJx+Q8aaOHe+xZ5kPr5cW0HVdhnJ
bvdbo8C2B3c2Fzmn0bUQOGSB/uN//KKtlI82r5aCcGDVcwO8Llef6gp+GDJaazhS
nqjblpYgtammqlsPtfEO77PjcEMh7TFC59uya0+6a9cDmbyNkyb6uRd1Xen+3nh8
gEzTiehumqiFfm4ewVpKv9oJtZExjUmj/pkwbTE4SGEFn1uU9pcRxMAj/hKhgzO2
ujZhzkC8X74nYmSKpARQltSMTf+6Ah25JYCRZMSFQ+w+9/SXgOhaQmjeFH++e5Ku
zXuOYENyT8ZwqrpYzEJA9t2Va8Utvh56dpEPphY/sXKyXnWNbPW6V6vVdgw5NLkZ
csqeeb7BBRihKUmYmwiO4FVNLTx6JivifRotX618wXhXpi6PrZkVYqfsPlxco9zy
oB+XCo1lTG1p021pnR800tHpLveUNugVN6Y74QHkh80SIWkcyReVUGnd8mW8AujK
yxuhmnjDbRiYXUvIqtCvwQLUFPOi5ilVtzen3lLRKJlKNXHz29y62ef7MPxhBHK0
QCwqJSlDfa60eN/HcNbE/4l8fYg4GmSDUzLITAQjovxMWQcd1mC9Ftbk1uwglfkb
cxGcio3TLfEpc1YH2dMrNLiZrNBcmH1b1JBGKqDT3g3+vS9TZc+pLFh/bmew7+hD
eini0RAxbl6JN7VMwOJYlh5sWwOOyZc1r3+bWj+oK2UkulAp2wFinod3wMGTARLR
78xmBSXb9DOtULkdmTA6aIpZnoGsBMhKpjlHJ7nZSFmTqTLiVWMMQUTjboqgLaoo
x0FUSlomRcziSW45YZIbLufcCUCUSBDlL0d2kA8jS70l4MRvdj4OYHxnJsxWHFvU
Ywfjem22HBDXSRTvhAZyYT3AGzBjHF2CO8ITAJ/H4NbHMTIOkDnNZ/tRIqvZxid7
shSvfS1FW/siTvQtFvYX3ZdjEY6J+M8YipS/HPgDrV54zJI+qGNrLxA0PgLs0a/Z
8RebHZoAie0B778YM/rdvYeUnhwhKoVlJ4L1fIK91TvE5cVWokgm/ZXX+W6DXJWT
Wm54DsjQU7j+chFaMlRqxaVH8WYr+GvL7gL7ijT4Kdu99PQTLmGOIETX4BvUVHq4
cQghMgy6k1c45Yi6zvQfurU1CuivqPL/MxGHUpEtt+O3B4O4P4LLQ8cU00tT+cQi
Axe1tYqxy8k+ENzZacapIqaNDQzykYYd6OsrddNsOmUpmqlsfvXSUn5mmYUVZdaL
VB8l2SOyEey4eyDDDZTm749T03nGDkVMUYMdUfsHkLsou2f2Li2HZrPM6d0BHmAJ
6rjtP7HhIl49CJk/X0P4Zt6XBVPh/rbMhcLiVfQ1tX5XYv7tuoyqHeGrLybBVML8
XxUeVUyLXTesgLqmnNmCVkeTwPtmfmmx1SadLMKnV/CvkqqXTgKfao5Ma+tkQnaR
LCXU6JCc4Ujr0Zco7IyrLiKNqQL8jJZBYn980OR7cPxnomt+LPXn+JYQwmwCa3cN
5TIDYKkITNRCnTJ5GKMPY7xm4R6SSZGgW//Ef2UF9HlgMpRHC7zvNpB1pIRd8dP+
PUnsg3ACqilI+GEBOXNN1HdwC/6jv0LMizpZJaSuYlPcbwmGv+tw/WXsAaIOTRfY
YFg50av3lWASHxUoQiEaJQYwtrWkVTFn30qlKhSVGRrH3NRGFNlHnr2tXWWFxRX4
8YMDxeGDTcTx0b5JArINPz5APtGf0z6VutPTSnwaF4CXNxGMn4RoVcjw+I3B9ZFG
h3sC2a461WqzmxHzNHQKKoGEb67igqxcBY8ftfM7dNFbyYyviCG8eSKuZKgAYSdC
IoE5zruWZ9JKjkN/7ROAGJ96a3CKUMoipbltb30k8B7sCVP/N+vGd8qMr6qjTMu3
7+P6xfpoPfsB04Yar3Kbc6aViEbwBATwy9WrhtFCu9D3qxYiDHaEjFn88G8LJioV
acTHzlNqQgL0al06c7oYaTAgGtTukp3XOvmHeOtla6Z2I28JLBi39XbfpMuIPVRG
gYetD63OdBP30XiJOl3I997xqtbAzQ5l5PWKuaXefqtl/WoPYDJWWoSLwWwNiGmI
ZDwyFHTgFFK8S0zBJa/IPYV7EwRHbw59A0CGNfKTpd2XNXCmv1SOqqzwquvcrPBc
RlgLzy79R2NwGSvQmYFMHokhj7SB4X/FYlGqXhcDIWv6d4jWqkjB3muK9wWsVdX0
pvhsBlLrQ7nLwoN92jl8EkY/R5fZn+Zb7rjLAa2oM+Py23/pGD6J+OkVK6rYVJT8
0MLADc5BIq8BufIhgLWw7jrYdj/1adO4SE41BhDYXy4sD39OIyIyY0ZeKuCW46DY
a/4N3cIWzRI014/fi+MxEOI1gDp1etqqMvHSdD85N+DzHqFj7YrUCAyuxpjPTU5A
D8UJX7rVVkINLrwJupu60jR2Ghck34XxgWxXwrD676lbFiBIGsiXwtQ183vJaiWA
HOVpwbNTxtquo2DnnbcY/nAPvRrk2mrGgfMdk5CDL2AvI00g650Y2cZUIL15ltR1
ziOkwn+26kL22yxjwTyyxs4/Y6yvl95OK4/QKKrESysEFLYFeLj1BbOEGP0hwP9W
CIGaDO/2dVhIY2jrt7iudARJ10dEoWxdmOBtX7A5nQuxcLrR98TED6nAlO6RjVPE
yQDDRZXSAmkerqkYuqtz8+w2gM4qCsm9z5iOD9CFSkg3uiYqyMyJyOqBACy3UsrE
TPABeBqPqqN7pJ+If+cKQSkKmsxnqv1UuSwBaGBUY6SyUBtKv58j6IgnQKesRc33
+4Po9n+AoCrO1I6qt7bG7HDGk1I6LoHKE2CXCB/IZn6mXc7JL2W0sxRkUHjsHVHK
gKiCADp/UvE++yef0D9LmSFO1rnD+lCT9oEcSpCru8bRU6dgOzD67vnnKW0t72pM
HTitQ8EQGCDWW3mtp0oiAOhBRFBoSlxO0FpMeB3ER7kRA5EVr8Tli2NE1UKBmDwU
mr4uvagv2RweTu1r7JOrtnjbCCqVIoLArl3k7UGijyVA4Hgl4sZfbiaS4o2zwRg9
UvMafKA+DJmma9A0KXKtpUVBFMl/8H01C6Cg3ridV70nxuN/NG0xsUOsojzdYDM9
TvanqkmuylpCnXbxnJLHIX1viK0Rh/dOUtzJq8rEgFKgpGClTO4QFCHbIIaXg5UM
d0MWjP6XonG65VmFyJ5DKrUwWNXsdoT8QLJltuAaGX32e+1XUyF/g1eXdT33Bw4E
nU95yCDvXSZla3nhcIFUl3Ga6FOT0IwDYglYleHuevTI0j2a6znwmaMU0FHAt+U7
Ok6SpVmXPFnik4j4npomsRbsnEV+0p7P608aUd67hSxabToE4QJfoGpLUqgfyyEE
rqP5tZpuVNzif4URbdn6hXwVJaEmC6jKVv2kWOMoPD7FmuaGTAA9nSEKes8DT3nO
SZAFTiVVHf5Sbnp8AxJ+ksfpHvUwyuMWO1aED2qHTqxLXJzf45waAJgRMH/YQ3ML
b8XMQzj0h6i8MhGMMcbgaJvYiwJ7WbCqRVoxIXnNBMdjhys7gFIVLispBcvdIXlu
MpXY2ZoHlcEE/F6rn3tCNHCNSy2RMqNxCxuXZEYw9603UyGcKG7HSEIxfoQuUn/2
mFFqzezdsXZAzaA3DN+yN3RTjjyQ32ALqPNJwp7Pdi2N78w6Nw6VJYt9JpZMSqgt
AcRCrlll1DyxivYsVqSadBL8yFNRMN6p7U6KNR7XCe1qnfdkHhkOavF+78FdR008
+BiHV0SIR6MMOqzRXoiptgp5IExkgtZOywTOy0yT2OytRhV4oyeUh+rjoKMsZkmw
Dn22dvUTidZEr6Tm942og8gOp8CdUFoJFFrmBWOEkkMSZZyMkS7MTnOgg6W5cH23
nOQrIAXNZSRo5DSHNR99Afiu1n8TIA1oMd+jhhVCK1GoPvRGgzuYeibX+SSdrV88
1KqCgPDidcvfQvXFttOKq30HCswG6cZXMsfYtYYh7iEtzhZAl9I1t5ycwJRGvUOS
fyiHHI1GnDeXxthyXP8tIB4vI/an4UQ0Q6iB53gPP0XDIWePognHZbwk1DtgqkIo
PMt15NIENNUYRbBfS+0NX0z2tSazohvzaRAdXfRl4uXVbAqsJaWfWlb/QFHQJxW4
Bv9P7i/p95ZwWq5LAHaqFPp3VAWsYKwoYCHVjKELr0cWreD+63GiDE5ZK046eJCE
2FVf7gJupVCq5/8kXZX8VORgokkONf6T4h5S3X91ZKw43w2lCUWPk2Jhe8iab0Ld
FI6+EOiJK5o84BAPnICys4ZYowe9ArOxlx1vN9M6UcBYeO6qxcy2KqkpxReNXT1b
Igcw3h/Uq18/ENuV8+NIPsnrgzg125nwmMcFwfZu5o+Rre90wnwcfC/ghl+XN3S4
Qpw/oKkqZ6E0gLAGCC68/4Ij4wRVrc6TCqfKfbvt45grU4fuwgrfdlLNsQVCuZGz
hjVigxUA7C7U0Nq2ZZeDFqNkZyBLg/zdKQAaz7l10I2fDs8TYXGxk4LJZtTX+puY
W0+f8N8BKaJiIICyIHOE9Xrd+u2lt79JI3xdzrcQ1Xvna63/uSTTnsjIaC6q1CF7
aE2wgBVMm82lT8lBOGOIdnVWKhgqQssgcNmvW6lHBTGKLzADaOUpfiyU21qSxYJs
BUZskyy7dLjoiEEbDkz66Mwo95guD3RDi/YkcKLaxJgYthHQYUylEKrCthQ72uSh
/o4415Dl7Q2wcyeFoWcnu0L4OA4lAs5BYDal90d5Gih/BaUv1a6rujhMPpyr0p2e
VcssWKt+UfF0TgnfDqnp90RkU9Ci9e+HZ/89L+6CQ8LPodvgJ+8ZOM/BH9cvY0BR
mDAYTMMp9gf2eQRqVXLwJDiIwHJ/svWHqAVWUXqctsTTvryWjhG1iwK5qsR8ubSB
0PKyiU/geuXoy6zvFmNE3ZQ/OTP3ycUCYoG3IDgpAhIgPe6n7huaRBH5cDUwrr+O
o7QyjwD/MsjznUEuLPnqjfQcwT1mhicJIqpR6M2pdo6Yqogr0XUeHUJFoktQk5NR
8vvA80SL2QsK9zq1jRp83SDSSfesAJJSN7X8Cr2QPL06evy1BQq0EuJViF2AkDmQ
Z7Oid09jSrqUE31eAiR1uXukpDOzpkAj97vz+adbNmrrwwFs4W1h3VCFkM7wI8Lk
RyZo+deBdWXB5JOlQT7PY7iG1KbCA0LeTe9KSLQNj0Jo3PcAvTQzESaCmzsiE2M8
uTjI+1Zb/hWXr5i4CZbO1SBzLeeJdXEAfznj5DgjMakosN9lT72AIQILCFiLvqwF
Mks6OabiacFuBQI8GHue2miYnufV65o5fx16vcNTVgEWfZ/EHzaMeH0FDdXigudA
x4vfIr/BrStDVO3Vpc4CB2LgrdnbrMp7iTTx6qjFQobhs0a/e5jDJ9kd0o9ydgFq
PNPbTwKXxH/JdECWbH/UHLA51jqYGs2gk5y6vAyPF7WaszLgnjvsFxEdFv7tqxv0
cOmoZQYVKkX48L67BEt6q3dl7uRXphehsbBOMiIVh0QS4FpthbmspviacVy45V+O
8BzBBTCgnr/tk0aBi/JepyfofjFwre3D/XFtE4BSy66xixMIy5EIZW/hfYuRc97Z
LJD9F7W2reEFNUvshcLXicRXQirMk4frajsnqhXFuw9hk96CrsL+E0b8EwtbDBeP
3UCHMbie2gp6fLZjNVNmLbIa5FcpmS0ov/8bYLLSmsDNiTs3hbibTjeknfFbgIsT
z35U1EPRqTEtLNOzb7OaCQ9/cy1f4e2OrS+f+watnQwgTPlkZJkDzgTvQAPugeLh
L8deNmybYsqfwjicXv94W1tL7ud3ssaPZjFzcDuLpirVVg3MUXqlFw/V9kxUt4u2
mcy63m2EanF+dv4woeyqW1BlG6CXjpv+Sj0aHKVuM7AnyrYBAWNeqRuWwKTSzU8j
2siObQJTERXDSEjOaFeEO6KOH2owuMqKJP/ItW5PrQ5po12DHykjgcEnrJ6k6AWc
03lOo0RXiyWaW+hbnPuMoU4GO1QLOw4MSBN/aKpfcT82m8EalInjiHPpGn2pDPK3
xxMbo9oIM/vF0lwv5M3DnobXIkcCGKQ6sa6465FwDyQt7E+K9OzyvWU9WbfYowgr
hjXiML9PmSV+EA8s3oAAAVctD0wRzTPX0WmFWblpbQgDjQtasJ8VTOY91w3GsYTh
soA/I1R0S1wfTiB/xcSk41wtlC1dq5TNY56OM/9C8StKO5lEK38LEpduXxpusNrh
KjtLsNiOnXZPObpQNLapo/cCafE3G8ZgULdMnQ4jiFv8ime6r1K2PXou1TVnikiR
gU5fCCas3/aU5i/ZGyzD8tjuEcy4Vc9lsyjG8DZkCM0hlqec+dHHyKLZphZG7qsP
AkWsLj9GSEP79sJFbDU2KKF3h7gCnv8QEoWuactrhiih4a8BxzSdIlXpsMHMYGGS
mlT6v3LJY6+l+lP6c5BPSVdGUiyGoZ85bWd9j4RPlnCB1HbFuE79GRDlCBiHkDuj
R7YisoBwo/smrwTdyzh0N5XA/rqY71g/OL89vUIK5cw928TmjdaQi7jVxpnndM10
lBK4g4u7nwJNq1hSHgeGoizLgP6gX6ph/q78/icmKMOV3N/3JvlICUr7faJzJwug
JOMiRwoduz/oEg/eShM5FutDRF5eFLGHptQFyUBWiv7okoBIyqyLS/yzxTFkOBRa
CpHMXqxPHJtG+tDiOFBtraiAloUuUhF/zMdztbJHk89HKmHRg5/YIGTwMZtdYWRB
fkJwfJ2MPS8mlnCObO1sxKGYwwIrVajQTeGIQ0ZIBX5fzzgg8oecbygDlw5BOXGK
KywH9DmDQP6PAt7n6Va6TRQsEiUDcV3zc/ZqFAi3TKsloucMYpWo0qf/YmRjqS5F
77gW4tHIaDeqHd2ge8Y7PSv7zBM5YlkxxSRoBYWFdNWKDv6Rbtjq7dJgnP/mdlQi
ZuhyE3X/3NazH++MyCUX6L6XtF8hFuPLq/NvzABnrT2W1wQyBOdxtdZrVSnGIARF
NhwJ0sPfUZZe0hgHdBpccJOhtnd7+iHoTrZbvmhNdsTh2p2+eVLer0XZ6/rEqM8X
12Va/H9as2UCaCz0o9ehjkgGaNRyYtUsCxuAm7Q2JsxtUDKoQYq9tS8o6hMmHkn9
RTXMaY7qDScB2xISo38H30H1tuEH+6Yh7RnZneMX9UskO9W9dpjswLksVQOca6kd
y86gbQAkkOQruQjSaC48yp7RQoz0SZC6dlLlUEov6QayaCv7qTeE6hzpmhuhHyik
vfo/0Gu61VgOCLOTaxBt5LX9elRuYpkr29j5nhATLMNtRf/ZoUBEatqTp75S3mH/
pR6Nj57Mk8kLEMRD8+qGj2dyfnWI0nO3fuMjbzLvWOd5Cy73OrSZbwfFAv6J6Zda
cpIry3OFIcIQs8sHmT+41lgW3s0PzwhnfZvs+8Vi65nPE5WavUfGKSDU8PgvH+My
iFqXP3rXxsn7+0HhNDbxpX/Dy5ZZKuNErFwg6Z1Xq/QMnQWsL5CXAMaxeEt9GpXH
xgyJdV+3Ui66b02ETD3qB47Z2pNsCPMORFWdxz1j/AdLA04UGXUzKS80mzO0Yfaf
Er2RrIhbi/M+1ZLJomfZQNgy9iCbpR8IYb+vCWt6r3Ar4+2a2iEObDgBuql0Kx5o
Sk9az/rvCU1p29lV5TBMv7U4j0NsrMbrGGOphWrwSLFz5CALHvbhZFiP9P276pjP
rwJs866WMMr19vFMDUgZ+h4rZADW1vAmKlr8JiN+T0hTnFQKr1uByHWE9qTXHtSO
MuLzZhud/IZXWs87Md/+veekYRVEmGRXtwMfE2rwreZmmrPQJisFveDm+S2gWdw8
W5PV8PmV7HpaNrDRFI1CvV+kHdLkkRKc8X0EGBrDeAZfkEJgCmVwLHJE/dzFdtnr
XpMyv7hRnSr3OoBUP5yRQaX7DomI6xPa5IuBSuv4AUVIvrV0x6P227fLOhGLQQF+
Auu3iDDYUgZjyRHEKmIKBACTy8FM2NqmD2dENNnfkhgTpeOt27kkwOYF6pVGzUX4
rifS7s3vm1CLpFVMpNCmAvt1cJ2p4sOpapaC9aX83Jsr3e1M8wWixQHRfNndrToT
/EqGUP2bYuMSHTO79Myf7SuQm0EQ6Uz+xneSiOxp/uY2cRinixrb7dTE9kPPG2Yp
H1gEWQBcbPdLqzQ7bBRxstn5maRJonsNaRLQ+x28SHzusdtF98NBXRSxSTs302KY
uWtFk4xnCcM7mWprgg/wKZ/2Arbx7J7bUah2C7s50ncgE1HI8xbnG470GzNUPJli
7XmDoRLX0WoC7l+BkfeOiAv0B89KI/KeGXjQ5aigfMSeG4N86lXdr/+hfqLsfI/m
bmeOr8HtAxgCLk2GSnFgsdBI/4QB/8s8GlKpu3sfmnZJx1ZYNZNmkMBfAFwge04e
T1/st7y2XuYJ4BHo53yufXkxsf6IF+DQo3/FRxEtBVsrjHHgYR6q/3e6LeIcweTk
1EXfC8WKrSX/kFIFyw5fXxBl6oc5UZrIu2GSMBAYeCUjGIByTK6Fj+dZzhLO/Vgf
Yj6VF/UK9HrmpNYxfdl/jqfXMhqRkZN4+z+IviK6rIrjj1EkKVjvMav9pOu6jkRG
jO0N59Qd5K8Ub58IFuAhQY9f8JImYoj2uxlxBDkVZgxzwP9PlKspYIkdaqNOvyr9
bMBGUeePXEfLrbJSDtGLNIACyc8IaqqrIw67OZP2Uda8KEHvwEaiQ6/sAW9vU2iB
64AETpRtsfCAEMRZhNzT0yfpSdXqL+TJQMsWJSULPhaB1Osf0W8f6Z2HDEAVQQ9/
x6UNAVbKvXtMGz4mdNjuqWdnRQU87lsV2UFvVasLaXsuDaNyOSbRNS7fKncDuBOq
/30gD6SfkwNoobQ4+7IELN7blM690lWFrtHmEtJxhCec3J9sDNzYmzo9WNfCb0Ey
H8z4keKSodtebJIpW44OHlN2TJc9OJpzN8jijj2mtfGmLivlBu8bazAqqI6IgBgM
JWFkRShCswI0fWPZ99+9u0d+cjC6kn4GBfcc8QmUoPGz0HR/jogWOuw+6lO4v17X
N1SrFhcRxznnWDieDg9xjojfF2f3vYuNyCcjyHraWjfVjvxHRANO4zOW+40flPy4
8XxDO2f2fnGUIZWiHh9sED55e+pFUglSj9CCu7Ssag3ujoPau5M6PqqvAe9VdOr1
Qlm6XU1XZIebZo5j+923aOUX7GqozO/F80PxA9W0mFhGvqPJmOmvLlMjIFzz9agD
sAl1SYVCs2qSB/Fc2O8iJOSBn69uwkBtQb4/a7yh4pGH6+i1wjl5NI0ayFk9r2Uw
gs3QiG9iJDIXO/6FHFS6IdyzTMe9+xCRhzqXq450w0bZTFvPsoe3nXBh1AOph3zF
LIwcAbdYYAMiQxsh3o/DRdZyB+ZSrKoHtmW6TFIEztP7KslwkfdwrDI9wJbDQYdQ
uOJj7v26BKU0YaDR+7JSK1DE+5typ1s6YEAywGcUrhHhb4L0yr5mwiS1Z6ck5GZP
KK5PrHyYaVdRDKUq4QAfDg8t18qM5R1qlpEWHKQpBKiKUkLNs/YnBo1oNbXIeNZx
IvY5M9ziSFKl2gwnbG370WNcOILhgp+iw4S9i4cWHuCu140ISU15ulY1WjcNMQ7l
N7FRLbwTQvQPYz2O68SPdi/iUCm96xqUi3IelAwQKdkj/uKwmK4bYYUyu2vG9uwc
KNJdCwpS4QMSmSiUXKHJ0cRHGuaH0rtZ9Rrh5AkfqZwV8yPAifIVh834iZ8CNTP0
1DO5wxb3oT5hsj596dcIvQojE1PInKRQ8w344bQ+k7UVkAcTRR4sa8BWfylWG6xX
ez/Li5WX1Fdr5+BXVx9msoyctDNuQ9cF8JzxVRgDKPpYW/VccbiteTIAgnDyrik0
4LbL2W+GnMjMJ2QCWeXuO0KodG34zk+zkIta5hb+awZN2BIgZp2pGbBYFiP1ri5g
FEA/rx5+6WFwLvDvDArWArLTu5ntFFTa+SdBJzsSvdqnrz3qHC4gtc06S7Gaka67
/uXxfZFNrY5s4gb2iv+aH7xlRcNjMjv2nhAWWdK4ZrDb2/WjHQOJ3fw1lK4wAtwB
7fQnEqHHfx+XOsAJD/zYYVtSw3kkk3sCyWAkD0C40sdJ50CiLl2wDiIU25cEvkpP
ir+/GpDlYRmL/PPv+wD/IhlIzUlKKGIiqNAqNJA9HcMxjEIln+KYF1K7FrJCPy/H
iCwO7yPCNHX6FL/H6Q8SZSpu4kx+sUREFyDACYoYITeYe+HXy4OPwdQ5UzZO1+HL
fHb4KzyDA2GunnaA8CMCxsvoUQQfgReqUyeNLz+JRY/7iWn1necJIvGCs49lRr3d
x8hHYAk7QMAPhqzIHJ0BT7vlmzpPlVUdjMMC4yRf++PSdq4W3lgoeWlxFXTZSrxZ
1S7nj250oAp3abtJ4LEH+XPAQAynNwpU9uGXYAdnVmPaKNKIDoZifKB7pH0/lWjR
lUvNaGjMFWI4KzADWv9IXoS8MXxTZ8br0y8ElgM9Cq7ElJIqYsQVS1nxtMtcfp3u
TJlC653VI7vg5OlgCGj/MUoe8mEk49DoiDvRKgsIrnAb5h5bXNOchQACXWA1TLkz
I0IJ6lymCXszaDdVfaoCTw4G5xe7UnSES4ibW+HssI9s7RKmvo1Jic8nXHRN0wo6
xlsK6v0xZZbBp1nWm/6kK0GnWuyAH7OPz9hjFntu3OLd97i4H+Ynxu7t/sl3woy0
uLhHSAbEB7tih62RHo24bPtzH8gALz42b0zUGbBn0U2Z6GVpq2hkP8foDHZ3TfWk
AvsOiLyq7tzroGHuSJ4IJy/CV679PFk4F2YKBepsYp86aTvh2WdkD52bZBxNOx4Z
TUqQskqNFHJrA0lzNNkuBLEEo2jm8zwONEOupAQ0a7+4BmiIIPZnfO4HDQmySBLF
VucAlKV1Uhf93D0X9Vuj7nG0q+sZKUJOfdAdZLyIYNGxnqfh4GEzXQwamgN83fsL
lwlYX8/KJUqbr0iCY4KemK8bSXrgWr+rCzRyOKJsssRbwiLT8qKr7xo0IczbmVeX
1Z8Zf+nFbsxcCMMUzVPiLUkfRdx/hw4cDxtIgmidw+jLw81o/muTwH818LisPCWM
T5iPMDiKUhrNPL8mOw+V9GDo+HQNsPwJ/WECcXjHnHY+/hzFPLUhqoUEWx+d5/3u
Avlz+V8H9OfKtBfhYf1RJ1fWADwk2bJyIP5OTu4Cv/uO1S8jIbmTaim0Xi4oPld3
azOt0Lc/K3RliM6PXSDwnpQ4lKI8lijo9Q00Av2E/Ca/EBkhzXd5IvpmPDjgoEC4
GsL7fb5ePGXeOPXbLUYi/RlHAHhGo7J+uqgoUvy1s498yrHBxay/unp5cDeduS42
tnrhCeIeTafRD8O8XNv6JQr1ndReeqVOq4OcEV4tZUCNGsGbAwAMTMzjmvukNWwW
JZNrk1cVRgmifGvi61wlFuFJ14+3E0BxCZ4wYzIQoLFut0hauDM8eYmdkwHMMHRJ
9zwMJm4EFQwasFtrCgSoh8UJTQ83qn0ht/pZ5nFLMDo2l6riHBG8rMqArPzOszYh
JsxJt0FbqKZ9EapDq75mizWbRBfn9qnQciRTrQ9vwaJgPC3iaDHvnsUFGfAfUzUn
GG8rSJsRT+pSvIKDgu+xKDnJSyzjUF8xMdk8BVsOmK1ZZyFWQAOu+8QgaYNWsgf1
IiQ6gtYXQzscBBq+he9rJKEW/T79ELEMx5XNnqRCsoIEJRxEkhHOa66vPo0U3sDc
3dy3Bfh9k0mjV6sPrGiv7eSq57HjUS7rPqcW2QKIQ/GvMgv0ieLTGY90+E4fJyy4
PYZfq24pbag9B6oijTP0htUUCEQg7Zq6YTO3GL9NKqkJzYoIZ+9DtunXRsliXA6y
0ILZi8Fgp1u+6GyLUdosKQGvoo6onYvPCAxwFq2mGKjWb67KHSXYWK3/H0L9tEr7
Tb1ROi+it8xizIasVuntNPTDYuNydnhkBAHaL8hdirvobZLNAu6NubzOd2zmq+pX
pwgfs3rijVE2eIfh43KQNpsq/7v7Aiqo1pFl05FCLfU2Tam38+TxFVoDQNfHYzYX
wC9XyRbglAUlZs3NvK6cYzi24a/6c0vD9AGEBHqqLdbQwxK02lnENuESW7ZichPU
YPPkmQPlx9aTk07+CgzC2oPVAOIJISLzEqCicGsxymoKtJ9+JYo11aIfNdDMdDsx
bHMQzyzXCpRbbdgjtCLMajDHtPUVConJetPpJoQDhATmPSENiet18OeRzH0AAkhs
yeYK4gr+NHOou/ij7fsfIrBN43s04esL2EuxZ8X0CGdc1sigXiiqgO2NfP4guu4/
3addg29bpCR1LhCFmtTuEWEyFzEiWmQaRtt0rP0HwUkbRvLXnvZI62Iw3LljSi/G
ktN0ht4gk3JnkSQd4gi2+shqVTiOGhSxCOXYIJL8ZDOQ+F6JAynefkdPaPEPGMka
b3CgGrUR3IKy5/ayx9q/cf44qPgbj4snUvHI8cDKFrVW82Ubnka5DByKU9UuKTOP
YauNOZdaSMIeLO1x8tVw9YGJhetIWzIXMxTDT+n1b5sPq0BwTVMFd1GKN4lCMuU6
H5913VunQNtGVz27BBkLtmOLpbamMCCyW3dmDn06tnMve56ekq2V7KLjGlZzj30v
3wrm+03GUKCwEKfPdE9ipHvIJwYUg5HInUb2VGlul8Jb2ZIaI9GD+Lfl/Pp+myu9
DAzdp5ji3KPCR7gyGz1M7VwuP2q/of7C/2wiEePwoyOfyFgJVIHiS/rD+M4THSpl
1S5vkAVNlYSkwvWbTEHRkQedZbPIVELw7Khowi3bb1KUM1sKgzQZ8z+qwuTqM1WK
/QYPZTcth7xVBjyh41Jj2gFO2663fxD747TWcdb3Nt/PVCl0IDALAAkEKKZGSIa1
BbueJrpGtE5VrVopbtAmkmL4/xPjOKfj5MIqM4UbLxVhqIMx/lvlhMvpJm+tGsaI
vtjMMi7IQ0lxUwgmN24DH7XvcIuQfq6+7jzOu0gG54S1jVUyZoq0deN9ECts51rm
AblqjMyViZpjjudaaHgY1heVXNEXyh1bxIt6MMyAWdEYF/D0xJ6CPe9hRta4xTwr
3ChwUc1Ov+DWWttfv++bF2W7BX0KnD5ZDxktQdiwxoMj9GTKHiXN+OkbNvnKEfmz
ZwbqwBwgShj67+asQx3vly88OFC5vjRkCDX3ITiXYl05xPNjKQ+endmtZleddHYU
OocRx2BianQAIAzaH+pl9F/7BQX+mCMIhVVY99k1fH2Ic32BhXCyMI165YBRlnK4
nVl3Y4TbeWYJ0HMLf/0KEjaDZEvB4rlWAiMWfFY/bcsyk6NRW6HZrXDC0k6BwE7n
8EqwM+btdGgo+ImFF6JLJR0OQFtnGLWe+YOzQ6oGicrijzsYWrY5plah9kgL4zK1
zhSni5umLWGZgmSZo5mt4GvesUF5pzvGCvg4OAvKBUpYuBspuNGwMyccup916lk7
JHS4gdrF1m0jX4azh8pPfn8IFtupNKdkY2z107gwxuW8D3Rc3gkXSVKWl6p4bLXA
L3P48FGj5Xp5gHhITsU9eCO1neA7kpI3F+Ha6GHLDY21ObXGB9L/yDxjFopY2iHa
uP6weax1fMMVdIyVQwKxVpGbCyBHScktWuv2dNrWGjTdok41RcJx9eoyfB7nrnxD
axVM/rWx4bSmiZRaXE83Jzz3ImGJuHtQjjwDANjhurvgk00BSlybl6rl0QIgldUS
PqCdywo1RkYRqdrCSTcqpTT2Lgk4SghpoleCEbgVbCwcmcPwVTXFf6N9UHdqPTBz
OVqLeK8EgMXmjP0aRJ03kPZQp+TjAe6n/KM7KCbT2vwMhJsY+bK1oPySkrpBQ+2Y
uoAcH83EwJ7w2PMWp8a9jDuyJM+K1zSJ0nuLFNKKiVaRRpJaoQI1lc+wjHCb4Rmy
t/MlGVh5uy6nPBuU+IQQi2bUDhbv8ie8Xtw5DiNG5n7qzJquxzw9Axy2aPJ5k/Bu
7J806jlzCXz8XpOuMqumccfNRmgMUkIxsjExlGf6MTIdx6/QmDtR4mkuhJpnbxY2
tYePDxOTf3OWpj/hJfc0EM9v6Ks8NDcTx8PXVL4ACoEgU7FD1aMrTU+FfM4M982y
BmnvRRyV5xEEib5vf7ZmGcqJeSTSzjLKIWpCqfKxX3DasotBMkVqGKZuihXGAN0E
b+nN40V2uuj9+eGVBKhp6rNeDoeP2RoB5eO3kH2/jDlMCFaBy2Rr3zSk4+wbUjXz
DUmK2xFFcqUHWQjSS9lBzevjXj2+h3qxKCq6vEwGdvgLdfb7YGa/1bXmAp9mm5B9
8V5dF03RhLaT4brdq5waS2JUzwIm8gkInVP7GLlnOsOakfF7G4t+p4I+zl+LuGwp
D1GOK1r6DQyuvAvu2MiB8o/1z2eu2+9wMmeLP6Qh7a6wZ60Eo5kdB64Z/IVsoCRY
mPATYrluek1E6nqo2LJN/dwuOXBytma5laJBXst9bhioZYCWzNEyM4UdS1F49KtM
49Xre0iiN9HtKb6/I90BcokzMTe2wWLDd2WXQoD82+gP8YBgwLBID1PkXK57OaKp
KSW4vyZ5lp4xaHJs++kMqd0VpDUJh7NNazYSeMb09lAirZa/n34nCoY9Y5gOiwvH
LdkOutfShHHJOvcqmu7Y/Nzu2Knoj8rTP+Ic81FhougY0IjdC91pd+23XrIYMHNe
obfsIJvN/Xt0/rBzi0915TP0rwx56oZXlJp2CFKLEJ3/gYwVdWTxrWSSW8Y70oC5
qwFZFulTEVeqdEDjHRLdNVzHGLy0fapbdkeXNnUIQ/bVSAXkKIuAAQrR6Xss0Wxf
Nzod+lAexrHcAM/KisFi58BVHcu3ewLScKDXspok1QnDXMW021u6wid6s52JecG2
IbJR1lEYUZpbIq3aP6tuikR23OPJo+5b40UprOvCSpdmSnPZLZJdg6MWXnnnhMTv
X9zRm3lYfTLVN9yBAAjawh06j2s53I6voQROxwTnSxzfaTocS3qNWzvWpuIgDzA1
fR/m650dOzIN6QBanwWHtdNrvIiA3tla+pnVPWMICAiX5JNesNw26/VKFZmgwq9C
e0B4GptSCtVj9Lti1XoFxogg5eN1dsn92rqxRieJnPmF7OSRTWHGGfPMlDiPJ33l
piI7S6SSjKoCiARUcXzYzvpre18nYQEkVjhXISpbYsJNsSjQrXgur2TTsNGuyEs3
aGMt8A5q4pgs2Do4K5tJNCZEjnBxHnTjqxTFta3XI20GRwdoHSjZfjXu94C7vJH3
RFUiq0EY74Klm6NW2AlQaxG6y9Sgtb+H0rnMhZWz1nFHYpSiMSDOzsKJlPuEBjVP
pHCQWl9pHbXCDws2kfC5QFxBgKk2mOWSydLBq4oDE8wkqg8wtrUzd+6SgscXrfiQ
5sGvNRQE72wGqvO4UBqO7Juigo0W6F6NxQ1MTqS+UYx9f+xXgyXmrxK8PlmpLGWA
Tbx0kfHwubUmMpyrNOvJB32EbCyD+pDty1oc1jbbQ41tgo6xQ7N0G6ayCbFCllWQ
T5l858bRXJuA/1eZXrG0uP0ucx7QgZ0Az0H2OgR78RWmV23BMxE8ap4s4QGSDrbZ
TiJBD+uXqUmJlFuwoco8nf0/RuGm9DdN3H51JicMtdqmSD9GjOSKG3fb1+tfTxk9
q+Tlxqu2BK/x/qee0eKFNNgw18A4Pnhwgl1gY4yHnDCDwHEJeELoduv6tHRO1DB3
H1Nx/ybiepUtFpGFqseHL12+zihYV9Qd+gTHH6Zn3YiKy/jMty+9QvAq++sl06I2
doZHn8bmph/UbNhK+j4rZA9EGK4GoVkYVI7/pgARZDHm+bo+g4BNUmH89MbpLw/w
4+Br4GC/jZ2xBv+ALA0cdv+KJj2QnQ4JGCxKaWSzyCWQSYB4IzVE2CMdzLTV4T2L
UQkXiKctzZBxcTOAj497BreUOZhP194IGUpR3QlKUSN/BWWb77Aio0F77yc/DwZR
9Tw+BE+xz/EwOzOCnE9ejl31QX3xUaI2/2o3WkPBCkL2nQwGI+FVJQiVJKO59O6y
W/rKANcwmd3QTlo/LAppFITHzY+QhX+1yqSN+AeF461lcWbucxWqnAPY49OHg2PT
RqD9o+dsx2YbTK0YdSj0TAXlKj4t7wlk7jbCtZ/eJ0zrk/iKtwwVPTcY5X1sjQEj
Qcu0BJStA+30w/xMvx42qiwaUFDqMdFekB/ypKbKwcwACKFq+Ig0EgMSPRgI9X6K
wCUT0YXltRh+toBu3lCVsI7OAwuzplK/ej3D5qsOxAUDxPo/TOCvF1xRGxTr60tn
+S5D5a+QxPNJQg4qNpUOPVPYx+8oa09VvylJCzqmwPnQI/kBL8LDaZWTGWEU7GNO
CTiPMwcWmEpmJYQhRA8LpFQTOfgpBoNw4FTrCPg7SgppfPnBw3CjNhQKzdV1ABtn
/u3K0y70Pro7zzOmzfjp0LSYFVKtKCAINYG5pxk0+RVVtrLNiQfrF7OECZkPrkJ2
Mqj69feiFG6SnpSmtFfbqqQPvh/Bsor9Cfs0CAGjgUCNGZPAkRGXtsdsJBi6xfSH
8PsZQ2xKqwZVwMxnFXzTs/QPAka9cFirJR3gbZBzL29GaJCbm4ytszlRnh3eeavZ
T1fsW8kItXtAevQgzcmw15yqlCCGVuYUxxGortLhyhthTFElDMsZTYB5ENbGG+em
z4B4aAU1YOm6xVcbSP/tEvAtXvvYpLAggk3qYcacw6dGgJyZVkTiZSIAtRpxmQ+m
a6BXbZhq578n9ECzO+gZqC+tl5Z92fLP8YE8YyU+jCHCEHp+AA/1TSmeFiqDqFeH
u/WodTckQaTr64mr+Zm1wgeOR6EQAEi55nm2RddQjPlMtC6+jZSZLlRSR9fmiwqc
JoxeMoKxX9ceq/JV5CaCQ7KDmrY7e7dj11mjHrEG4BeqXOn+DSa1BEDhAfePuGff
L4joc8JEguNks+wmgGOe/ungbPfnAdxMVwrmE/0s4if/TBMUMz9fv4wzXhr3nxgo
yKjxBSzmukQ1tLZNozAm+EgAeFCycXuUYfkJMeL0nbyZjKeJvxF/us44Q27wQkPc
wXlvlY0Um/f87pFLjqqblti5ZUHiYZnQ694mOHOEqvs7gke+9cKlQGh9UgUBxPxp
4Cuzd+XrgtNXeR8ETGM4vRsZK3Xm/dXyfGlGo9K80Pi11Gq1CeVgfEpMjFzHcQ1c
Cyg2zdi+qnabBi2d42Kqe9QMqjFedLZ+3L3wt0DhabMPvL5oJu/Wpe9hwYOj3tgz
5MWwxQL/3iEHuxQ6mchami8mykRMsSBfQ5ZFtJ5sAlBrBpezyR7EqqV5V177CvO2
fv76+r0fNZIuFSd4hUX+6Wx8KSCrkALbXfziyBNRLw6ijeM5ghMxHG/ZGqp1VeWN
JfIXf9qgvJvAFzDbJXyFRg457tbxvX1GCI/YLat9rggJgTNpaIduLhScSZbT2SJV
y7QZTj3inCA36PAEIBKNNiyxfBWVe/ENL/spSOQwVc0f4GrKenGn2MgU4SuqC5g2
asqVgetugoROhEdqfzyCW+ph/Njko3hhvWjggrKeHwTNRtJlhhG3AUOOtU9hEtf4
iKuCLbxLXiWDYZfDfZQ8I01Zfx8UwX1u5hHdSspjWebGBl3+71GI6Vek3xEsBS7t
lVOJmbHStvS9ZfFDvx2g84/yilYvuhl1RfvXYwdNwUQkEQ7IefUKTD/AV3gwN9iN
qYSMlCZiFb2nZOYylkxk/eXKWpwgkmlhx3EQLkdvl57GNUN9DDMNKTUAhRTmllrM
H066QFTUiB0ql6h33IjFqC96aS6JtmdybpyN8P9qcAb6VE+JCNo5CcLAi0mrvU2/
cdO2HXIFo53IwkFnLDNjd8Bj9kg1QrjOsf05zvGYl9CdHAKJ4xfWjuVsrCpwgAWh
56FiBMyejlZmtBG6Dpf6r+uydeL4v0+cN8fCmzMXbzmX6SlYXy63a5yICPN1bw2N
w2qKn2rSh6EY/yR8k6xp7HUhBiKjN60wF8wCcFRTBC88s05geYy0mxV8AkGMmyYv
gP4XyVDl9AcX/a782k83T0bsgAmazjqyJKPFFap5vJFzi6jhbIc3Pe5GTCPUf5R4
Fts1SUTjrfczVNO+xSWy85fcBYKR0TcFBaGpjIttahlHmFlRCgERvn2e8ug2gs5+
rsRIGokUxSWOqqgLlwY8BJ6MQqCfuE+W47y0qhHb5GDH3datFDIixxfIr/yJUeUR
i5j4SbOjCmIqs6Pi+ygq14/rZ6nNKj9vrm5NCzldSOh+dFsbIBCfY6JXcF9o3BmX
Ybl33lJZ+7U8JfDummzfNmPFXdQG+/3c/fhbicCLzEKS2kJr2K5zWTea4uVkjqF7
yLie0QDXF7tp0q4isn81/AOqePHcwlrxdXlz9FbcGAqf5E8XeqMPR+h0Qh8eXYX2
joPgQt59o2WhlpcyWTEOAiyGvT3gOlCy89Ydr4wbhYbwbVx9G6dY6D/mCUeJPdYx
ftG/SfP91D+6GdliQ/KIrSMPb+qUDHEpHRpB095z0H5lG0J4TrOY9IPT8Eg/tHKK
LneKyKkk1Bzb198Tsyy0kG9Nxs7EXLeOhtK+WZ5X9QIPCkobX6VBN/+Kkyv/W/63
qoVFAR4ynyGLT5B5y2cCZd06ZjAZWVLmNWDmoWw6/9s2bkO9saLFEbU6iAuZvOT5
nW4czAEGbX8qhLe4CbIcpMrqUJYP4hbK5L/SOGfxTAuXtfWT7Yl6dWrRWgQxycdN
egvOIXYEkq9F+Tz6UDFGh1yZI0Zhety6VQdVNc6ORoKcWbNwvCVXJ+moh1nTFYzt
Pi9S0Zdlfacd6Jl7HZT10XxPZmVuKccHx57B+OLg4QZ2lD/Ut0lrrMDCGDuufrsB
Kxbpt7aTkIv0/MpQnwX3yBnYI70WnyewELL8E6IKcMvMjWrc8bw4iGXnDJ3bQlEE
9CNfBXRLJSYL4mTMJ7owUXcg4tNB0DakLWX+hJS2lvMPTf4lxzcNpGIg7JHfWEfv
KdrkstXM1wGkMZPAlg9npUgWga3Ou9SzAEo/PZJzaf0EOqV54OJnG4iy4rgxbl7C
82GOc5ZCKfZXpitrbgpWMw+17hjOI+vI16XCykhkfIdtfAQ6MFqz23XyQrojh+JC
eJYgebH3ijxtEcSkdrNp18XFL6YekbBgViAfdDejzcqSHWHJ0fjdrVayTR2Fkf3y
7Wlon/IMGcfY3rhi3eizO9yCE8qad2e1C1QwWf/JPpHVYs4fRbbLf0Kdx25Ydazo
M9Ftlubqmo4aDQIG3nxAdrvayjFK9li7vSQKztzbm6lGJtjn7Bq4yE4b39dkiwFb
gTWuOOL9o9xq+qmrGz0NkSWxZKvvY9XkLi9nCPx3x2o+LKMUkJ4pwr9MJsBgBEcF
6RTM3uLuV1Oo/1aF5ed3hG++K4Uk2vT8PmjRKat0gT1gUzSv1QPKTsaRALgMeYhD
fHVCYFCDYMJpj6ItWCcIUPLP7lXOxGZtcC8wFsSmxl4+CVtXXEN8N1nUOsvtzbAA
OuMIBY+7aGya7azwgtsu9AR+l6E00yZNF+mVn7TbOwvlqqTLi6MaX/J112KGr3T3
2Pbj9/OhaH4CUscvnt/wrKbRBF6R2c7m3B0RZF5rkfNx2C7lOI58oeyhjedS/1D2
JThfz1iy+ri/GfxJGh1W2ANw730yzyOGd3+kHNEJbRBdGngCn4QekagnAgUnNDhF
agtD+Z62s3jKH8Zegk+fEFIPfdxGdlxTZJFqUCWocqxkSm282IstvDRxLs2OGjjl
+bI1QeMtotGIziV49dhKW+TUlGWEw4LCFBJyvWaaxz8U3Aho/RvcrnrN5xJXlEBm
pjTYNkAaTSRwiEtp/ggGChNzI8wS9kQadEF6UMQ+iVpd14R7McjgX9TpXtQKHglA
PhV1pneaa9KrMWWmSmGn8isXDJH/avTL4KUF6VLrDmjIy46kfpO/7Ul+1eGesAxe
x70RretKO7rqZaYiARQUxt5i+pDGOTFHcbiK+UwGHfbIXOcnotzwbMXzMpBUzaQF
BgKpSXYT+XzVunQCRO/esJrI92frp34AhDrMTX9oKb2/CZ1/iS77T8mlYyuenFkB
ZZXY+SuWjrxkqUpAto6DjImqayB6tkKpZspS6Efl/t79ufeJHi6H0dCZ/2R7EibB
eWJBia0WVMYhO0jsuzt7gy/b0oca9FaQwSz8mVdO4yBkyk18RTbd5F7WqzWWZw5C
sD292ghkDC7mDUeDEobavd29fbqmsBUQARTW9eIpHfA79kQiHMeCaXhgOPDY8I+R
//V2vLBaNzVI+ZOfb9OpJcQNMA1bsXxmowL+e0vD4hqGKy0uPzTaYTl4MVzYI6RX
U4jHC/MxWn5XvgfOfPbaoxon29sL/UgM52CuwcOCMza6Qgv/Qo17QHo6a8EFg84g
yPwlEXfCG/zdZQZMnZINA/RcykLmpH6PZOKGX7VD/egnopEVIIGYrCXcGGk+W43x
6+m+MQc0lZwFpaXXZtmYLeZzcobp4tcUwRDB/oGBMQyQOPuRwYk8j3x38ZbUaPs3
SxcqaIB2E8SOI+BBi5OQT0OSxk3ecaTv7z8pff0E+BUArzuis5k2GiJq0ugQtzkm
/sfruTPS0ie0aNdaNISl5b+Q58U6QqJF9vuJ97hscKyN5wAw43hgl8Xb2R2mhaXn
UOuWerhj0gQBB2D3kK/XbwQswspjD3WdQNQLAZ13vcSBcSnPxPsF91msI2Hp5vB8
6YnNKed9rox48dBDXD7/muCYxOqoQQoJd5XPaqkmGNOMLZyBRwkKW4+wf93HkObM
5C2P9hOGlOsZK8WXiKeEom2WoiXBpf06uUTIE7PZw+uXZb8X7rjCXXmkm+z9LE6i
4u9S51MLaPGZfcvGyJ/xS9pXsMsB0bmLdmSSXVEqvr47sJ+Ubp5jsPE6hIk8oK2/
hacKPhwmZUo5kQA3ExojbS2uCa56gKAaS2c92XJS6Mc/Tbp7+JOAYJwB0+2wEJop
Lo70RVy2/DFfBxsqdWYOghocKodjcaC4pE8bpl1esbwGEXzkYTI+khyrn4K7j3OO
KLefFerD02lyT2Pr9dsbZBtJ/0W0/K429FeqLwaryCh5y6CDKgELax9tEpPkNy7w
hB3AeIM/CeKfUZb0VlLHEOAESyv4RFUMFwxTW9CAzA/+AzzlTwSBTY9rhKQT3P/i
FQejMzZYTiXkpDzJFZJseguwfUf59c40Hf5jeM7wOs4oJ5vonEzLlmfygFbYoavf
7g6pDu7jkyQFkmCfmXyvRsMp3kSodf0TzlG9KmevGMvsc4osVDH5Him9mGxZGzQO
OEolZ77Y0w7xbpwDR/ob44zxbCzM0y8ZgQR4HcCgEyKPXfo43WNx66gIyFwS3tNr
qb2L5bAyOyVbAAYaikx3W/MtLu0agmixUhHtLQI5tJFGVMiWl46IOnmLgCS4RRk1
Xjnz3IYUVJ9469Dcnc7P4DGSg/YoxOJM7yW36lphtISB24acCDlekQk7v52DII1j
dlGQWf6vs5KjhFoa6NFNotwjyrVnnNut4BEbsQllsTL86k8s5jsJr/UJlABsDDha
Wy7XQDfGshJsUJs8F7J59+ZA9p/TvwXq6u+GA4aXmCySwmi1ZEYvp1xwr1NFZxir
gfo6Yt5hORxPoAqg4BrRoOduKTRBxGy7JBeH70TUKqGx8m/4XPQqaTSI9CPsxOX6
MqHfbwTsdfetnTsQY1HBw4DUaTR6VnQu69MS+15vTZ87+1H46WRP4zwAtEfKceHK
Gz8x0fsEjE8c0m92/foac6oZMyt7X7ACVek4o48uNVReOiZSWeki5ZVBDIoVg83I
eQL+42bHb/Ug6G6W0hk8BMREqszSMtJmhIY+dbkEmx0fgccLOt3N9A2xYD4Qw2fE
aTds0L4QEhdCzpgSKglrG0wq6zh7dqGAFxZO0z5PVqXRxgEdSlHr+D1yXi+6q3Vx
RgjUsCv/NkHe6U6G98XCS5Zll87aQxbqDqA760xlMKz3ZBNs4rQKCNekH8AB63p2
sUHXTC3npq76l/lMEpBfmpfpTUwO1T6yw5F9Oz0N0Y8njmTNN5m+rk9yOn0v9zMS
7gwGkH+YRfvXik4Wwq1Cra6ia5YCbUGaFhcjFKgUgTipVzzOR6osnwddta8oY50N
FJivNb3eFUE+km+XU4zxOeYfYYrQKpl9L/ivUVwKod+Kdl7CxFwEbJFtD7SPyTNQ
vXN4IOimozHirMCzz6j1bzbs1DUzAXMGbszWVWtG8QRKX/14QRUsawcej4b8cFdD
Mp9YZN/TulC6qVzUlJ06OE2rIb1nsfSIFMmC69JI+EijqAY/1tpbRfTVmbbjt1EC
ZSwFTyTj7RvyA2c67BBB7n1P0YYrwLJcw0NXHR7SkGqZyV9qSSUc37VSN/j1GznZ
5RXj2v+8arm6YniMUuswg7lmgYEB6OObxWMVH19XcmpC9Wm3BvA+9y5neESNHkZr
zOK500n8FcGRa/DvtD2XmVohtnldOiHx9y2mHqVoNo7+oDpQIHyDFMmdTFLdWVw6
7DQoUWXnZQJ848kdwuL1h1Ht3HS2n1VuBz6QfZwWsUNZwgJj8LvF46nErEo0uDJo
FgtA64R5cwEQGxTaaxKkSjP82cTmMEZMZgNyvd/EdykDcfxRYKP5SGVlE2iKfSw8
2noh0ZA/Ztv9jXfoJShTu/Xovh8Psu0XrJdILL1P5SuHvKKcMpZTXQwHbyc1Rvm9
MCjhRZir2ZlUvKnPM/ID/GGHN/qPCDKApfLpjBt1hc6YhV+UiYq+7gEOuRPrErKF
dM2JYI60vZg5KiTienzHxUhhN8b4WPfDOwQqKjQ1GRXK/demoo1YWnhgqtsMkB6T
zB1U5Mopx2zIja1Jv/4nygAwYezqmZngukjZVHkJtpEoA8W/8th4jZcSEqAT3A4N
uNeL0N/jakqyZI/oy6W3MYA/rQay5tjm9iSMIQeS6xUr4oGZvUFoAVKWWjMR+yhh
6Nk1zKlNmiZ5e1etf12QXaZrDsq0GPOeO/hG9XyYBp9gqtzdz8Ow17/bS8WzK76g
PffwodfuupFj9ngv6xghbHpJ8zoDbfoUCIfH2oYCudIjDy+wUhQtWoRjTWKBlqjZ
IK7RMjqXYgjHWI70r9ANJa9q4wW7eQi1fdUgKkk0KEoGv9CgaMWmFzZ7VSOkFHwA
Y7y9ipcJpSAZuYOzFtSJvT0H41LMZkWEgeCZARmat8oLr5snlQhGG73rY3ad7j6f
gf2sXOquTjKcy6op096bmTOmf2+7J6npu+v6s+N92I15I06zHs9Zfk4ovxexnOo/
CFUVdQ54r/ofMwNX8Ja27Bl6fNH4AdmNDKX85E9FxRSGnfrRONdkMZaAyfOWYYy+
25qdD/tQvPKZtk5Vx8NPQtqSe0fI/Ny8KjXzTxX9FaCmCrBylu0xPL5jPUnRXiCH
PWYSK2MWesgNeHScQ4FAGj2PpmvWY3auZussrMmnRnIGlTdpEROF0Ux9bnYrTl8q
RBUx+dIEIp6CCeZCXDfpzsLKcv/zOVa17H+5WpKq+WhbkuAwyb9eVB6ckMmgdXiY
xv1zfPsOBFSHeBdDl2/leErbmXSJrZy3EnbtM9UpdnYznBHFxdIyby0yk+GSTtpC
vclf7+9v1mRuvAR2vISrzdr2PJmB99K7oar8GJTaUeHjwztAMVV6zPWb2GRN7GiE
w+FCIpVc4RXHKOvhfyiDhqAR4nJ9jppMryGQVWC9RqkKdPq3A58IIdtKWs/0Jqd+
ueMQ9b3//+Nut9LjpaCx5FgzaU5wxKe1snDSJg3TINMYtzuIc/uhNAc3kbpGVKYT
NiLW0qPL32Zlu6LP1oE42yso/OCEZ7EXoper3iaKeGC2P5sPGDeQdBVUrPrVaZ4h
2jihrwHLZ8k7F0ePm9PxARk1fIaqnYzk7dIAYQ7aviunHvDeEkbc6VcZyPDe2iWe
6qp6dDJLtkA0sjk3PEOsFJ1Jiyy82/GYdK6MlE6HgEfXjeO13YorLt84EBXY41oP
s2MbhLQ7uUYb+EFZ/4Na9MKE7KwDEFFyGn0EpcYpFGe1FqcU7fpzdcLMTGd+FlJu
RU/2VJKusGdy/5wLj0IVgGH22StFj1c8hGO0n+jCNofKIJmOA6U+d0Onbsp0hoe1
+ezDUiN+on5gVc3+2glZUHbNq8eyk+GG5/ZgBPLm1Y7Dp757U18NA8JsQ2VlPlAJ
Kw0A63s4Za3PWPgRLy2p7Iu9Aord85wX/yRjqrZ8vRJ3tOMhXQSui/7+6nticviN
tt2xo5nZ7w0TgPX2gjblIQ/M5e5ht11WhwvPj/LLPAfmq28Dmra/E5d2CeYyDI6E
NKmnbKzxpMCD7fQB4h0/bZJ6Y4xSSw79omlhQC0Y+45K4iqfXmObUX1mwGvdkg95
mSqE3RWhktRxmsiXvYkJ++Cyf2Te1iJrs1na9wHcZ/KKXuXa1O+hH1DVK+rm/afk
ixmbgeFp+wx3/Gz8Fb/xr+F1cWjGrcj3ryk6feex0VahARSv2eqC1/mDcZkvkJHw
F0v3cGjsElVkV8me34naxqHJtqJuX1th7YSGkq3bWux6z0ou09FHSUc4aBlc9ZQu
fX04Yv+l3qayWuHG0PM6tvhj9ao8kC/v01r7mCcpoSAErSQAqZLzmtR5zo2kOdOw
lwoJ1QCjgghoxd8tPO037GGSRPmhAfDx9UAeSLhTDpzCuK4z80LiQxs97Qesaqko
snOAgWMiZeR++Ah4+Fxw3AianINq0mYr1JveRtIaRRvt1nO8f7LlM0jxE40GtguD
Kz6jI9lx/S6w++K/O2y8rxzdi/AhSHhmJ7e59/OJdSiV2tAN3ShvqFcNM31InHWy
RTVQPFBUcIgO380lqjvIHrX2fwba3XHx5Q0JIWkWPPp1rddBU0ec8vH2nm0rasbu
civKr/MJFTX0kosLHwDylGRHBJcWOag4sOS1chbIYSUnyZcbRdYJvMuuQniJcHH7
SXEkEPTRAxDVC1IY2AaiFYwdZWmdeFLcne0TXitbZ2ZzU0xp38B2WeurrtgAaP5j
zkk8jSF6zMzPx7wxNfYp3Hpipm7FicBQkwkP3hFRX9qjUGqd4C7juvAcSyGn1HQp
f+t6uUDZD88B2YM9/XY9/VTgAI9mrBcvpGqJZyoHrzG+IH6XVMzTOvqPtUSg/TXY
WHkuA/6igi4uCi7VA3DQ0wQwLm4EWPbOxzF8EkF0PxbRYBJnZaNc1NhSPI47a1Pn
/UvTuYePKVWnLRyF/RniQlzwBhVOrZrinrCtsw1/NaiRyHLB/3xAjcU6oXTnLn6e
QapDd/jbXBOrKwmf+YwuXhDqOHAHMR4huL3G6VLDwcjM/l7cN0b7ilIDkd7gcA6Q
6Gcm3s2Kx4BJxFsUT2U0hEl4AQ6TNVIDiNAB2LRDfg670ISsuWeTVEyGm7jXg+as
UNIAIZkHy7cU81Zhrq5NyJBBIbXxYtUj7T/wnmJSfaw7TlXbz/dk2YwqTFsOtqsA
Z9W2Ye2srUIA8zNfeqY/ngcgFKP4mAMBtmj77N23T+ZrvGbI2ZFQZ4UxCoEPSMfV
tAEiXfsiux+yiBkXeTwuelBlfRjzZts8wR22Da/wILdf/hj5maOH3a6IvYy/xEbK
pvEM73kg+GqXRjTYYox7eYsBOQReS1iwx7Gh9YpOPMNxDZzpw4lqvBPxVzzfYZtJ
etY1MlGNRgw42SX+2HVdmPIs8abOxAnP16D77LfbPL2fzXR+uqFmExa9X72dUzaC
EoUyfSwRuUjGwvIXaaKZLajpYt0en0sN/Nehh+zhbUGFZmYDm3TZLxM6tTOtQ9tn
3evX91oMf+CI8wyGdcbfskZ0a5HGzHt02e61WJMwCXKz8ZQyEIxZiI5afrtOw0Ip
9VwrKXXczZFnzrxQmD5DaVCGSANMsPD6CMFBJxYYIQTKIFvY6s4oasGT+v78gfEU
pK3Xfy59BjeeK4PYW/eBm+y/FBSka3lX6qiBv1OlJQOZ5nQ72+4eydBbWI0lSSNt
CoDdC4dsKYstpaNoy+XmoAXwvKn35BXvcYyfoLROvJxqeeCii0+m5e3SQNxoA/l8
Rafg9MuuyP2MyWe8ccNe5ZGgauhSTgSWdcv9nm4XHcHWci5i4CIlprQHEQsrv3Pw
e7/U+6GAu1aa5UZplOl+5vT2Mcm1d4zv6pfhbQLRU8f23/T5h29F6C1Zp5i1oDBq
nSXa7gEaApEFSVr4j3rurv/f6RGA1P9rj96gqA6Tgoz4JbJD1kb9XWWYmQ+jfu19
iSobERYHwS3zcSGBDVn1C1e+1tDG38PyxeJe897BDKxvuGoAmNqu5eM1ILRZpAXE
tI6gHco4US1kh4p67uCi2lNqXEOjmHJVd0Tft2a+rGIJkT9EICzLF6+/USjHhyur
CFoN22iykXb8bl3OzfNa+tGYbWyKmGTqj42qhR0TLWTxWtLLnIora27kDgijWe9C
cEzykFtquJsVvQT74KUE0hz6VELRQkuU9DCqV4dIT2h6GsdBue8vDk+QTYJMFMRa
lG+h2GCmpjuHpHl8RTSZjnjZtFHuZyzxVxIVx9/Ay+op+EvdpeGaRQer+FR2Ieh4
1t0yG5OPHkhXQxj9SZEpCFstIhaMwkue/w58bV1exNV5teOfDX0X/7L2fm8gI6JF
N1loUxSUPjuymc0Bmwzfm56eig9xrUaYhGzrfaOCYd3CQ2dEvOVV+rY/BWtkoDXJ
riJ35y0UldlEbYtnOzi+ytjuYStEQEghaJF0vRRl8Mn2aTdt3Lg7+xULh00Rqn+1
m99k38Zp54821mQiusGML3xqe5N+/srjQQQSYJlm9zfDnuCyRkwx7ZR2UchUbrcI
TRgJg7S9XhHyC5F/7c/Bkp2/t6CioSqrCko2Qzci4ri3RbEi1vVaXzRyRrCHaKmH
Xsj0+QaBPwIQYY+8OxmyemMydB3uHITdV8X+cPdnyfA7EeMzUT/PIxA8MFmr4bK/
pZ09lpqdOIuD7/QWTv6+1mbJUbnTwC1NOWoOV/CM7jU7dYPfnm9EJNASfBdS/Quk
p3Yu9FeX/SYv5PfaIrsGI82SY2DrRZyRO8xnnhhRLMUVCn04ps0q2LNQmYJ5xsUd
RSN+h9E/urKRCcEcXhVqBtBpthD+2C5PD/uJXuCMd+sa4VI1ewKvjfUH3v9/RdM4
PJF4FTFMJ3jsLYUXN6mDAbnzVb9M8GPXR+imo8tsR/yZ3J+yYApYHsqh7scF1tBx
ou+0pln7A+OMU2mYcqIFCLBFcIoHWYJo0hcFAlX3RnO1o2MA42RkMuC6co3VeAgZ
VgzyswM2kx94Pb7UnkzPoCIfSsNQj+6x7voKWzXSm6z018LQhEfA2g2YUAZ04Z2s
EvicByFbp4pfF9dK5zjeY1hLXG/8f/R1eC5NKecu2szAx3qM3DMfaQ/laYl+IyHm
M28dPwS7Ejm0NA8Ba0bf1BD3XhndaP5tECpYdLa2At6Yxh48HmWdRBHbda7nLbEH
vkg1kMUmeyUEOatqVDBMTv9GlyiSfpIsmrHpP+YhxbT73DkdLbTzvF4g8SXsn8C+
M3/YGdWXJ2zXMNGcXdFwXkkALLSuYXylMKWOQvRpABFhqBfL4VkU8AVKrzBmCHlz
/z3vNH6jne4WLai0f6ftq21Hst72vlZm+izFRzgd+tRNoon2ZSXSJxnCiAiThUiw
Vii5ROgXQjZjRJso0SGyxwbhb0T2JF1Dp+Ae3lQ3FlurTpIR/zlCtGq4CRAEZEpj
p7QVOd8/Sp3K5YDqXCpBXDNXvLAgm3fUu77LGsC+ZKrZBdlqhd44VpZXn+cNJ/mv
+0KaMY/RN8yqJBLFLa4I01O2y4K4UphH1lA7WsEtB3GpHBwXK7TlwgF9D9ZEL73J
j3M9LcwM2HmFLVxManPlePmWXOvJBud8XAIOyeNU/jaLRz1WMNVBoGHeThHbZkJz
sK4CEzp1uup2TqIlSzZO9Y6Hbqz+txwloTQZ/xgLl2+/1HYH9tRN/OD/4qhwKBAA
WKqAuYWzvuE03+YDbkFznKVZs71kvmGqP6O0/kn/H9Xzf3ic5ur2///oINGNgD1I
QbxQ/hJDzFwL6xUG/HSJEQmWMoBQrSJz1XGhZSBsKr7KGDn2tY3yTHlfJ0E/opHO
QpYdTn1Bp8YU7L/mN80t/MZqD9p43ORpfO+j0YEwGxSBOSM2ZMnzx4QhYuftZ2h6
WZ7RehT7qDHYSl4Apv1NzbxvT21iYdFG/Nl39V1DO+sF3CHqzV7ityeNrM01UKhF
7vhgTRYcW4z2ymVCce6sP9nLa9J8cJ+aNtqQHjcO/qUHTuzvBOtiZnp9gWVUULUt
YeJPnl1bCgk0uq94PQvaMaJykv4gPzeVgD1szRRt3rUbLu/JzKYdT4qOjxlCBsAQ
OYLrXI0SXHt2woUlTieiWKlfvHl90vXPxQvjDel7yX93u8uS8toYJ5GIEebp2PDu
UJ3SVoIwexIlWCZpR+IlBDrgB4+jpt4cpt4c7X3HmqhsUZ004eufkuvqWm1XmJEL
IwgF9KpWDnitsOMQSK1Oq1uAD0lMIug8/PO/aIXX0q1/9clhZL76x0afjOjNADXm
q/RhYIW3Lrj/03iyhga/F+5qBdCbkvARdkClFJm/BEdfHGw9sL24cxeoxW32QDn8
jdowToEZSJQHCplh8LpcrRB/p9CDPZxV0WoeAzln17P61J6F43abSSiaLr+PobAx
Rz0UEewI5pdUDYK/h4iPQD/oFOd1ot8Ta85u88Hbs0W/g5j53KyG3WOqlMNEAFuw
Uzfjxn26tRDabP9pk9o0ou7ZGYUqXyGT8fYxZWzYg5PcBrfCq5NZ5+vV47f/4q1i
tJyZ7XubxAyZobbnvzF5oTJaakJZVO94a9Nya5x28Tdv7kRIlHiejYi2u/oXMVFu
pHd/PciYNB643uJ5hT/9Lt/Gonzw104JVy43Dslo7IWkVKiOus8hfn3ZXGaWLRNK
4WRS6zFGKMXeWCn5Cbkne8e/HBnhhmxOTph3huj/6w4Tnt/SEDvQVMVCX4D1WSah
2q+0HgOcqtHWj0OQQlcT0q1ndt3rRVz7oRLM2EXAzfhqdiCsQH51c34hXdRseMZ3
yfVcINh7QGeprGU1yEBa6wVAbtfR3/woJT7WqvI6w7rXsFTpnoIj2StqLNpMLjh0
/Ke+f3Pg0nWWz22Kvw/4JbY17MN4PwfSzwguxaZYpuiX+1lW3fDIt1DFLvwvg/xU
E0I4AEoJKcpxFKvjJuPA8bS6CXLfbCn3JehhPQus/VdoyrzXf5MSoeWebP6hzU6+
D2emwysbBM1y4q2fLogr359CMha8iW95SAKQGOTA6Vl3ncA1YY6ZcC/d4OKHmAwj
RQGpGbORxtfwv1pkWwbxfncRbPGp2AXqX9561eQ9bsNawi7P9BHu6a/iA2HupJsp
wbCCKGt4/RQseCKfShLqMpffPH0LjpW2doCPIDKpEPZg7E0FQTf3iSt+iQkcIETV
IWVn+j1dt3UGnln9g8Klh7PWC6ycsIJtzyMWVMSLEd3vRH0YqSUn2pcTeB3O9pfm
vwXqlaG20ZhXDKxCQ2GzuEDUxaxOa9Mo17la9fjywm3Rhe2PyX/H7k821r4aASP+
Ob2e1Qnc6efQEGfEG4r9ALq8P25crRBmq4Hi/j+hVh1T0PsyIGEo+r3GCXhxd9Yn
Ildh4lbrw0B61r9FXYeMp/TeN6Q9SmzB000ZXymsZw53ccslYNBZhQF70+hh5jkf
97j81S0Ap0Gmm8GrrF5nH0MZe0SgYMZJf8jRAeQl28IeIoDhumLnMMiugLLL/jgx
JvfC3I9wTi/KoCmFVoFMRMLi0FQGR5v0Ylp9LbOinxRRqnWhGPwKu5Uq9llcyx7F
XCUmN9NYVQEs51E7Ert8wv++F+79Fsrd07pcpWvcd1JQG2sp3aQA3sWO5/Q/2pV/
8bA3wB9038PK7suwRWlGJJZhbibVP44WpJA25r3q57q8zH26gOJiHXGVESgOFXUL
r2wyIZH2TZqUjerlBPuG/B/sWRFN1m+e1EE87I6fVemn6V2fjeNVcP0W9bx09K/q
WOS22ZT1ZnxKzVUR1kQVeaM4Gc6ZZwhFNT0QCAAcoXksXXZjUBMELb3jsAgdBFBg
r3hJQbeKzay4SgT5EIXIypO4EB9TcoVlxvPhwymLchsGXPfAtmHH9APLA6OI2lnP
jME4Q3letGC+5rYLqgmb3O33CdMAT7EVSmNLYVH/Wzdr1TidDN9f+sCtZQO0aOBo
nDyjZTg6S4SLSzilgfyvtvJ0S7NpvwWImeRxtuh+nJankOxtVX9YxyPzOxs1NtzQ
rVzINO9ICl0e8kfZsz8LSYPfYun+dKAehNrI5s8MEO/5NPq2QJ2ikxOUuSU584ak
NSJw5Wc7Q5i6f8xPK5aP6Gm2VnVcaj0tyOHuZleLuh/ujpHDEoQR1Zb/O8ICjRnx
lVda1SMI62ovob/UcTSX1D0LnTy+biVBq7jUjfFJGAggYBNdOnuoInFuLePmuxgA
uuhGj56wrzeW9FhqGYj02BmJMpDA9tI0gxVrm3wD9qu8nhEaWSvqi26SgRKk9s7m
U7QfiwrmBvN3wOTNiDqz4yYvOSwfEIqbtj842bQHBoD2PcpPCSQGK9dFpyQrZfjg
CD/StPzPXyBUFjEYOu0DjpuKGdCCiYFsj5emqj9vrfbb1ifLuGMpnRBZc35V41rX
xzR0FlhVjyurJT26+qMmyW5/HKnlUsqmZfxGTNyJcXp9/ivPl2dTLmYm7tMpUCIu
jVwq6nZ1VRUQ4ujQoipyNOeQWDSm8KmadF4IgGGm6QIyG/YoltMPO8QGfRBJ2bpx
+iw8bFKGmnmw/Gf0ifTqSwSDNhVL3gfOJ+iVyOzQrpnuKjhWY8GGOU6fJyvmgz5T
93h/qxRccpxCtm+IFt71YlUGApd1xEybLN8CkBCQpAkPBnI5muZEHhYJ14aI1UX4
J6B/uZ73WQQ8poIdRAVxDQtUp1LkX+s1NGekkOHhv9bESMz8gsPDVFdPcXuvEYLF
tQK6zgq/Y67nn2xY01Xb3K7hP8CFeiUNeWJfpCml395/uXgQqLyyyjqa6oWaYxv7
52xZSVNpIBqqu5HcpkJ4EFZJ4k/kSBHauBmCJm0f3wvhoZYthmoNL6Pt9gFcuCYF
e2vK8Kso6yaLpdlnkh4+k8BJyOAl6i9Azhcxara4UFay0Xk7LfEB0Pl6w97nShpk
qJzBwMljfhZrg4jOEh6fGK9LBYypwu6KRuF/WwkLQrRni2Rw0vR8H/nBQXUGNXwp
8Ni+N/tpj41X/UD1CYHW/RsX5fdNvJaP9tl/hqxCkSjNY5z+wmqy6Py1ciQhwc+s
40EJS6CH+y9ZI3CeRYyaZCc2A4hGdP00MLua5qcb0XQ/NuB22w4clYZvudCKMD7t
FzSJz+CVMzE2ay37VynFeRySk8+h6VRzDbEFXi3rNCoe2+7Pe+HBuNec9H/hEBk4
3CViyQRV6KQXhpJpOrO+KDN+X4Gcnr9xs3QsoM6pA8sQ5n7+PARVwWf+dPbg/hZp
VjHD/6m8/ywcclH026vBMFDdig8VoBca/uEMKfx163W4Rn/zq7j1m8r4gMtJi/Nu
J2CuhzJ3oQbqBu9OfuXHyN+DHncoXvE0YSEAHizl3E1pu1r6iGu8tnofTqj4cGam
88elfny165lufRm9n0XWh1wIF2qNbOQNevV6WAdmMgny7L0JZ3Z33H68nC9BRdQ7
bHC1fW4PD3KUN+4QJ24//nfQ8LlBMFpMC3ripfCVpq9zGG0b1MNYwMgPl0wX3Q6U
LNWaojHX99Eymdz7u9q9IHAJKN/bA3eMbIH7WSyxp+kJriMFi3/QnEuGbFFzSNJp
9lsai+H5YkFa6+Pgyct7sp7ovp/qGG4mQz4L/lw6VWsKMdBX9KFhE5ekpgT5JdWl
VCTkKS5xu15AjIr7wg6sowRjPcSzr+YbKU/nihSAN8J/Ixi8y+TRZnkQypAqhYLh
jjVfWOR4C6i5qRsT23MzzKKZBM6VTdxh0I6Av75bpuyt8FEsNyPcJXZWUDhhnn8D
qCcSgcn7/fD+Zr3O7yCCkXe+YHo3TWsoTAz+XWaFLzpESJQ4xinsfsr9C4V7h0ny
UU558tlfByzny4c9sAnV+cBQXUlA51KBxMWGYH+s/OmwgPg++Xlw6Ntj8WcS0gjQ
lO++N37pjN/v8xqi+NzAO0h1xKEDEz8HDj8dwfx3RlYpCzQSzA50FNeuv7yFX/QP
nsC4ifq2WT25RkXV6nw/cwG23aYBxrvWFktZcMCw/41XSu80VdyDtS3q4OpQTfsr
eMnlTcw9QwEFWvrBR913Vq+jcr24kGYIVetHM10PA5fYtM4XHvos2uoii3dsG4xc
mt2fNmWSNQ2FKCuWoKLPCZunVVxJJ1gSu06hcdkjIESVX6nNFSdgxSfi3vW3GyVu
5JPxqd4Jx7U3SZOt2Whm1OuPRdltV1iViVzwcNxLTJX7S+NDWYZlwb6727QRpIWl
h07Ox4lxPBGkUUTF6r0Ro01GGaC14/Olr1hqn148BpXrKnI0KlutOAfX8hg1xIo7
ABiT3/bn0Gu6t6Gm/PBs8UjMGz9kFn+BPn62jWJ+lDK4Cjh9gIs5ttQfVXmd2G9N
9XIAfU4M1oBAtt6+64TcQj+rrdlNlQRVCmTJ9wKnQuLln6ZcRtNAD2nugdqxxR6+
lQ9+pfAM2qz1KXNdvaYKf8qtGXEtedS6XDiLeaGrUXLQXGeps8gcVrYLzoSXxx12
bjB7lpaCfs50jHR3WrLlsGd6y1HsHIhhiuxrzfkON4GTItt97WfyUDSs67BognXd
0fw10yQ0Zn4xRv6FR8Q6jt9msiR3HV71vcu4JK6A5dVDsTcxeVEyOgt1+khFVgFT
M0CDIOTP9mIGNyik6e1ORwYIGj3HY/K7sFVVZ9Iid66wHAfZUU2EjJV42p0taNVT
ucpU+uY92w+UnOKS7xX5rzh/MXQxlpJdFBEjYFm0PtEgPGKcx8c5colvZv02468/
+6jn5MTksHCS9GkOpMjAa/BX31wxu79m8eCXvNFT70DMIT7EcSSlHoXJv+tTTkaI
OyAC3UTIQ8lSrkdPNSEa7t4W8jMfSFIzGn94i3+F1U8padKwn6jld+7PSlfQe7zR
36IQuhnJWknfli6gMaIsJI3PBJEQsWLFUdufADeQAJm+H414NplYfLUA1zUGkGKf
ZeQVIwMFhYiTP5vv98ONC1DoVDsLGBClnxHxP5f6l9KyVk3dqu9od/tSjOzgTPIs
N5S4azt7gzy2H3AznRe4XmxDORFXJiQB+EGbJy3TLwQ7bD4d4MbMgvB/2ulUUiWw
rMXQiOJUUnMo1icu3QOC+MsIOUo4vhflQPyVXMIs3qad2PFBXY4yRP4tJ+5IrT1r
6sJFNQIWGUHoUzg0yq30mJ+NPRgvMR51/QclT3jCaUhBkCmFJ8ZuCX+AtB8/AQaS
Pkbybx4R3xryvki1cVV1DE3AxFRV5lVUvQLeQvCfAbAsyTerqvfE0p6CLppCdb/A
8Bql3nKIwa3UKxWf5cJPvJyIYHQxXaTy1cCqQzvDhmxM+FH0kDX7DsWjQxZoPXFB
q0AYW1RxQ3USBYmNT4GQTnlFfSRxgYwlnqjJfY5xNA86byS5okgxZAEIa8AGJZf4
+oqgwdAj8NGKckFLmLn5G5HOQhy5XfVdHlcwg+nT3cK5p5cul2AsHxb4GtaQ5d/X
5yEQHrRCii/D62KHrx42+gRqKhaKFh0/rCMnPiRXxkKtAoU7kGWT4PZT0nI6Hxsk
MgYYmJvMVRJst52LCLkVY14NXIr421modOGdkjQ/zJ55DL/KitO2STR887STSIPj
1RbgE8A9fYwMzrZTtk8M3YpeeE4ZwtMK8NxbceYoVaXvdPhpja7dDRtUUi+Kwnu/
DApOxluXRQEpwkr9IxUsqEDwg+D3HKKfdwRol1EqxIMqWzh0pno715sH3lxC6g1h
z4jXcG9vC2WNc89m5imWKA5RXoaEskfqZD+bOHFmpEuz4zpQO21dOaHqxRz3KvNS
NwXeWzgPWKMxOtBRrn8R/xt4ukrblprLbtb4DE/L7Gjm44kUwlzzzK59EDTREQ5W
Zg4UMkqdnvkpdSHy6L0kj73/6xh1RLHA8sI/3C/iigkDoK11bBJsbEiYp4TaGmeI
WNYtTIOqJBaCb7Z3Mwy1JdOi2/mR/jvGH/PwjNgNtMhh9BZOqAgqBhH3i9PCI9di
MU+vz57Aj7XcnvD1Z+0B87aTEAq6hgbJxXix8D5S0qXQtSbGWo0G0ctTl1vOdbZw
hDtw+RSq9NeQARRSi271ns0Y8/CB/csUEOWexsGtk0cmWbHxZLHo56vKZOxWMhcx
CL27iI5sRPCyvRJzVnYvx8ukMkS9Lsaxw9Z0hdON/Zt/v4ffhQ7tZc8/B7CGd+c2
aLYoCAnMA7i1njC61bNCYLu9a9b6Tz9Lx4caTvuCZQwtYulhJg6aQXoFm9nlRG96
TXfAl1O2ESkiMK8hYI9SvLMlibp3txWoGwCJAnEouTPkoWQCZhcLmTu89VdD71uA
FD4BOWKNRSL2373yyS9pRp8xy4MIDqRCKN3GL+YCnCQ7Tf7k5XjPdbjUxJhXcoxf
xSVt1Zaom7uvYv4cVoA3RMfFz7HY72HqoWIF++ASG5wUd/EJVSRWsEB/mU0Y78YD
AqH3ss6kOhFVMIEVX8+9Ycv9GVS/YwRehvs3zf0LC7nJKnmMFXaEsO/qRj7+M5+N
1j4fSNRFFbpUq515QAz/+9dElLpVXDZSb0196ytmSByLfYJklXupAo05eqUwqECG
zb/avy48UaTK9mPQHBONlOOzX8HSp5e7YGYPaxpE/jq0BWD5pZnU8UA5mKKShB3q
9NOxTN7dPi9KbCZWLj34MKrWc9IVfyNcoIi9pGqMZuQlZ1Eb6YTJhgPbg/TD/aHn
pieEMnuA/kXCcOeH5apQjIdHzO9OtY/MsfqnnkEy/i0SWThgcDuoXttAQTSDyTkJ
45ICAxdjqg6VwNsEvlCdGnRPm06gL9r89K9WwykqmYpTfV4wD5hVTVBqLwdKqD2d
AsqMfBveRkoLqf2hHNPS2VYBtCqht6/+LzF3E+tc6NBp6jSIJjJd+ZsKYY6gqFTd
4PQX0ss9pc93gZ34lgfGfDFBplegxG145cbOz+yA4BESFsRKPO7PZCmzzHsngZv2
CdK3f/uAlckSwvU6feOakHfXPwCn99y4fwEV0R7jI2sr5TZfI3qE4nJOj8mthFH+
Zu8cpf4oPSYniFpbh7vnJqjAlaIwIzBupwuBBlR5gdfDIiwCkXZnZTLTTsIr6Kd4
ZVOehMPMAo3GbvtAti+Q9D3UJRO4C05J2rekuqPLRFEytYCi6oJcT5kXEhgERHIV
7cXdFkti1OACpoRbU6mNrCtAz5E8OdGpbJydYQnwuvZ8LYnf8ZxHTOJTy1HB1aIW
AMITIqDckfiCBCz2HtA8Pt719x77+6Mkkh0tDNGJUl3AGlNum4Drn0jeBhSdKVqg
d+Y/u5/kEaTM2DqGmsmdmh0L5r2g7m5h5VC2br92Z/EIFLd7CX94QZumbnD7VeTr
bXwPbiTTrUrTTnJMsEdNesy7ac1S5fYOPfWr4jFvUWfpFmhhSM9pKbzKO9r80vFn
I5eJmTLADwuyuEYnIFKoVES57ik7XApOgS8YYOdYyU4H+jDyP19ZNt7YJRkxKdEo
4ueQ+RNTl+uvtM1bdmBaJ25+VqpXsL9Br0ZqPHOT9GkLqOB3cHpaDu5mcttoHz6Z
G6CTORL1TvyyhfNF3iM2XbmC7XjOF8Vc7OfGpEGXv715SMQSjq+NIYf7p6d2Udj8
vabZ0WObF8OaCE0k1t/nwoKyvF8XasSnBfbokCw98dR84u5pgooAKiIdNGFNqS61
iJ6MHWEAran9ClPlTZrxMHfDuIPQ/mZ25PZzivg4+2nMt8DYILadSpWCTIod+8PK
hDvNUyRvMCeYTFO+EIkWvw7iNgim562CiZT2/GDC5bTPU0LJSw94bSZF9JwVM0uS
SdPS9Zm2WBEd8CZ2FgALz0/TO0Rd7T1lTkdstk46Eu5dA+f4WT7epPsJtaeyiaeK
NSLrRRPII2BJh8Bh/397by5Dh2Bew0ytTzMm3Sq1UaI6Gokq6jUhJHoi8bcgKR/g
GKKhuknsHjjzOdt3tDAH1JjvclZ/GibOTp8jxWx/WCh3qblRe91PVBkR2BfR53lI
R1d90luzXaL/SqnOsQteJiTKjTw5PweJvUXaRwv7pJGi8F2VEFItRptZZg3usuZ/
jbyeCvLs32D0KvrWkgiU0QvMcWEnzg/8eGxNFE2KRVCQbQn9LmT58qTNr5SnRKiz
c0orDm98iOpxgd/Pnz/905d81/xKS79ywnzFQQX0tZJrhT5RnVqe/X8qWfU0+8Cy
DWnHflAXrOz9sYZejNQfV8Z+24Iyx1QkzHLhpLaEXLOqcOelysXI4r/wPujx7k+n
N/1U9vLRaHjTTH4ODjfxjVPwPmevuCYVZi5RQeVIvltnoLoRIf5u0sV7KmVG0CJS
7T2odHAYBmC/iaD3lmrGaN9HAQGHATGlQW5k1JbYunLlfdzEt+SihvAn+ri2OfNc
oxIx+8dmNv7os6cfKpqSCPRfmlhxm3UX9kzwYHRZZ80Iw2KIXQQ7NOgUMk/4kV4/
Ne9LlFDr+EvFXs+RwbCQP5Bs6ASbJKVg1qvPe+g/lnoGHa2iCypGlD6RIiV0ZExQ
yj8RSsnrc9num9PFsBJqROa/3ylytS4Sn+wpDK/oZJFap0yZDpwgquMd/NnQWoOh
kEBO5B1uBWnE9EZuybwaMmIQs/mZmVR5YZ8DkK/+iSE+KHP3uiruI75qPGYo70UG
H2jiUVO7+dlC1XVEixn29rfUA2ZdkzxFT8rlhC2WoC1BduopgLQHMzurXcJD9gIi
xkQfCcmH5gdlphRMkz8vqlK9o3Uc8mVPpR6nqF6duwdDbbT564Yk+bvlJRfMXPwy
8Z9CIVza+3z2zL6O4e5i8nCUlxD9jwf5aBVZR+zO5Tnn8kuI4KYfZlskmModIZ7A
OtLysMuoDM9v7AxpPvKFQHWHX3nwp1nsldmH+c4QS9BZn3eHNff1+CuKXFn1shOD
U+eQeIZCtPaUHYzzrvJAFoYcDJdYAwVJsZmubMD4PR2Opu07C5o+mMJRIp6QxqV8
rEW9HqtJZvs1wA0PcSeCtyXKwI0cPyu14dJMMdOoftlDEYB8lZzzxWvq2zJnNp34
aDZocu9TXA3tGTkJ01MNQGmUEGM932h+YrfzjrFdAQ+6x3ALD95I5R5rcjDvXwsw
PM0Xztdr6Z2dddP6fl8ui3NSRf+YxSPU+O96WEWuFJcBwKPlAdeGhvf9XD+aU9QG
VeAuJlD2DBHLmfABRBPuWWhssDPMyFdTp1PY4AahxPQb15BCP/k89uBMqrv/8LtW
a1vsDAouo2I5zLWIDn7Qg4HEPee/1qc+eWhoDTtrloMy3BNocTziFvryt/7s+/oh
NqYdWKX0d7US2TsFYRzzgW9CsaYH0Atf1VQHK2CCn/4jc0bTsJcXzMuBK/ZyUoB2
HOPAnjaEeGrgC0jqduySUQ+TEt7nlpYV/jomnEXrOjtUJ1Jc77Av6w1WL+snIq6Y
1YvUrXzBHF6ic9S1QSMBDY77dCVaZ4AaWiwQft2PPEfTSCVuRSJilqqlQ+9CoddZ
0TlYQOheOHHHxb8lIgAjlEn8j6LPPOkOsDWv4vAaCAA3q4kQ+H6AY1yMbn0NiMqI
7gbIfyoWIV/38DRwI/1zOZhi0QN9GHozkpDbBBq5+yROh4WSH2hz4CU4OVKFGUTb
auZ7+U0mjjjWuUZ1LzwJsQ5gzrWnDPvsm6RFOlATNegE4BX8y+AgzEmgC8N/yUPV
j6Su14sfapUe8JTahtpZ2JBjbvIhWLYpkP4m7dbdtDXtQnpqtpENwoIBCnMJ53y5
xv8A2LcaeyHgOR/FD04zFzJvbaikDGajcrTTV3HCE7uWqBCgz15yam4ithQ/fKdx
3obZEpeWQBr5l2GHAvja9nYEQIu0ji9hXWDCOiHnKzeOAANApe4WOVXNuSfcUiK7
tLRoiQ74IjwHKVN2jz5gxhazEnGhi+O79w+3aylPlJ0cqPGE1Vkc63fvA4FIxCbR
MfsuuaMION/rCfP8HYeBv4BwlNzy7IxRslKA7fhpm4jfttuc4NQROhKzXq9gw4Cu
0gJTqitHyXpczoot33+tOja9KrsmteALD4VZQ4xIMwTRXcxLKfnc2I2QpS7ZN5ZB
x5V7/Tb/d3uznV9PdZk/FvllotL75r8SVPCFIPOhHRGu58RibK/iEtSa4du93372
ZY1XfGd4888lDSlmaCSwp2Zyx7wvNGmYBJ5EnDOA8JDySYMk52y2DTa+AWs3cZ0v
HBVnXGv/lszSMRjiFLV4lyWe/WkEu8KKr1bMmugO1S5O6Ogy5XceHGIWEQbvFlBE
uIlo5jUo9mBx8BoR3tiWPTL6zoXxN6jPJ4MgQ/PimHoGaXdXv6weX+UY8ACwxTFG
HuPW4oO1tJWpf7uxETnQKLzKtsOHif+Ks2eEWnPcgH+W3//7mH1ZvnbIWzRvxuUX
ctPUi5J6qwDqnePlQKqxm/dEXCm6dgZXeZxIRsI+S4H90jNCt0Z6dyD1Tn8tYw0g
qMni/wjOKNFIsELqPla3mSRBSYDrbL/fxIDJ5Ppi/9WDM2bXgf/oWBspMOyleslo
oI2dXg8rwtUa5hvzV9gSxltTXmJzLaWSj7cXYq2AFwxBndY3seYxcZc2Hh2FxmXc
ugCv/i/R5XnWfkH3EpbmrlD1OCpHfX0rSw8FxTwOKHt5aF57IZ4bnD1VtjXdXTRO
ODfV8zNbgaLrA9NpSTi+/CWt/X/31oAYRSwWFiuLvAgu7a92EEtbEYYx/IMJkDRA
ulH2odsexusQp4YfS/QfhYaGxgFx7hxs6xV9KxPwZNWilCQHMiWWOdu+dDvsydFa
xi6dgq2J4VVoz36p75NaiwkTXwFMfGyeBWXkbyscDrrrnnoc1s4016YJ3eOj3tg2
X1KgiRtWeb3TRQpP77250UIP2vUPKaq9zKSNgegCidJne9DZAZuKAd8vKFFjllm9
6Fvs64KCAUtXhpZxcbdTCGT78KhO8Y6V57HYbd6bQwyfTDIUVPtFFmkBzaCvvCXb
BhDPqvi2fdkLEXbS+/O3MolZR0BZtJstZnsDB/lrzYYkFdoUtnFB9B5pbr25Jn3X
gtsW1KVZbE524sNedeXy/I+7m3A9I/jiWHIlqkxYLycwtQdiyQCL8fL1q//rqUV2
bqZWv7aUspxhv65LwNIkHn1/H/plKiKNLe/jdpIItN63th0TTAb5khdV2OSDg7iJ
OeXVZG7XFU0pQWuJdUDwtxr625E7T8KKAbqCZNH6AtA79B+nQqKVJpuC4CEeX6bm
UJLAECOcF+PyeOt/0ieiRvVdmY7rb+tO9BxP3qILKzK9sg5ANoTXjQk2iYBlOa6R
39C+D0qLxts0rh9ZIfFVO6ElLXDEj1wF/at+00g/WuztwCg1FWIfjpZuEhw2vEjv
Me1G0HEJ7lclcNSQbgHHCDkOK633MTPoR6LR2Dlpu3nBoZnonY0Y4jOojmHD+1BF
g+Kfh9JDr/IgAJOxVGTHQvt/EvRiinGlPTLUaL3Exi9ODyIc+F3j0++EvcO5maMK
MxsQt8GLDGQ8UYHXtHHkiViZJ7OFh4cc41hhVq8hQtdDHmziNKg+EwFRYgagKXxf
Y9sdEDlLZSsNAwuv8IT8LJ/NBQh7Clt9pzuN400wOXvdFflEThilk0+VX6v6xeAF
rhUGOxaYVCyI34L6b3S7jNV8uJtlKxGXnZT9LD9wszRJiiZVbinY6cxE4FnkM4WB
/5+tM/15Pg5yq67+XkxYGDRmSYfzs9H0dHAJim/ls5AAYGpuwNKl5lbfYhrAT9i0
jFxLPP3axcUB/M+K1C0dgTSMr0AvjRFB4/euiOGMb1A0FzR6xUJrCDlHLuJFKUmQ
6FEZvtyd/Br2PzTSA2Uq7RlhfvGfOUNth7zHA2YX9DiSioQfrAO2pzXlMpbSHVGI
oRdyYTY78mxwgEPZ6iET4mhd5IVgd0MN5RBWqIlpiOzCR5hNUEp0VV8nB5Ezg0rD
ApkWuWJO7ZcLgd8/5wuz6EvAfJHSOfmmO5ubbIuY/gezEEWAnukkSq8bvj5ycREq
wORl+5PdPAUCRLYknlyWYFoWUmARGsua4DlDxa9VRNMZidLuKcFpczG3mOmNRp1q
mbI3Vnfc5xj6XHYfhDvkgVbQdIsNMFYMzwgoUoAwQ54TZah3ENkv07DLa95LizyQ
TzcRAGjhxL6tf+E5Pv2Lp+S+sz1rp5LJobFacLDIX1tlCgYOtuN/FmOJIdcIkZRC
9Ib3B7obu1BB5GATD5uDMez/8W+g3eHCtE7ZjKYbHLlMTghuYGjZphyZQSuvTTLw
bLOTnxErqenHMFdRZA/YxXBvLKxGKLQAwLH3LpTZmZRY1aJoisJ20lQ5wK9KV6Tl
iknxOrnfwhZ6CvGoCa000hUMhn0SFTcvuP4KoQNArZoc9FkFgoSXmnhrEG0FtkDP
sy0h5J7XpZ7cEJUtFwIALLwsBobLkKzBuiS2Zo7E9t6LA2O+0A69gcq10LkAcygW
qosM1xzdSH1mu2nNE24vKGMw236+Zovl3abLC5kwP6QpQxesoCGsB9k+co9sjRRP
CUVGsmzKIVHLlHKxNZzMy3pIMTeI14TEE0oROndvJgE3IGg1qhcDf3E97XIWuRb5
RkLDg/rAxj8D8/Quxn0LAVNVTQWGu1ez73tPiSwvbK+luizIVZs2wiqHG4k/Mb4a
UMOdxAkAdMNOPj7ETzfXgiRoxopfF/rVc4niCdh7ohzNtR+RdjxZ657L+Flyt2re
ArNfG+sltb+tsZeDa+PV8LWSOF6SPT08/L7Pj8G7RLTeYavmTViB1gUHtGDagcL5
mmRH1gQiA/T3+VIvGE4Yytv4SvShH1uXynFt25eRbCZJ7sgmoAFwIlWql5Iua0iX
ar4dj5fvDlC676hJAuDfv0yPGPnqjUPQRjO+ZPQ4PIZJheq0Gy93P4FwgDwh+paO
wSf7Rx3AmqMQRSz+/yv3VoD8XXgU0mqBoSdhZ8aqEEbgO/HUoE5orwjc3hHwcS2F
edtPrOmDbuj4HWguk9dFjmZYHuwqTdQ4YgO/kdLqCyBo+0lEbwsqrKP1d4Pol+vF
KdHyEDXZfIAWI5nUjbOTbMpw2MjGHCNfb++VvmNAW84h0dZqh4a9+wjuyFGeqj9O
oq9SWn3kJteOojw5Kegoh4vgfkqOs7ly8mDs0SDI1Dt7LUSDPOR3lDU2wB+wl5/0
644pX/kBwK2n8r1ikf/+tobZeH2YbHWG12H87ujPYdYwABQT5gmAUR3Vj9G/Kllt
Az9QoaaboTOhyoD3fPOZNlBkR8PL2gv5yh0zzbVVk46sZngtBc4KlRffVrjkCgqx
YIeacobJ9B/BpMucuni2Pkc7eplf64bQyy23Fm9yXW6594or3oMxPBZjCCJ7VjEX
5AM8yH+Dhdj2T3+UXyzRX761ptidHE3TZFVV4zQsnBINfbi2bzAsvLVr+asAfTAg
Gi5vsk5ew2Va0bVy8fue32sV95iJ33jEq0th8soYNQuffMFMsyD7HEo9Hpn46c7k
r6IYV6OFp41WEcZN+Z3wuj0BDx2qAsJ+zGEqDNSc5vFckB954eQo9HVM+SewtNgN
YkHzladOcDJCuUJA24+vX/ZLnqszTNQsWHTEPKXwoU3hCjEXZlu1WvQkrpqy0LA0
xCXlbruk25rOrdbcnN/IU9R6KnC711k3UvcWtnrsIeTvIh3ML1XIvrXk1NwX0EYR
++bAaYsUyiKjTDlFg1jlemRBVu1rQbYHco0hJwM36y9VeKq3YrKw82WcMKkHvxl7
S9R4yIPQRCkP/y5yHSLWYaxzns/ywwh/ap64P1CEMnHyWPOx9RtKcERDl8lMmGwk
ARkLtB+58JjK1RtcMye0YjwLuI4kXsmAlay42Fzp2JCntF5rlws0vDXBtSmvqWcf
n+sA52Uwnb+/tD2koUKz29HtHyLHBwgh2AlVhkWPV5JPl5+UPXy5LJDrtQHfSFnN
yaWgBN01/omeIFOJlydqv11VNdTmVVKl5sLhkGg/8PZyPSTUMUjxIDQoJ232nm6Z
bD6IFtrl2Ic1T6H7eV6tcEt46dIji0ZBNN6MIB+5tRC9Gk9Nd4Qi/3tOH1MtoRSW
OzsHthDekLJzTO7cOE5+6xCT6pkAmRxh4QlmjCbP7LaMUOMNdF1scXrYynzsErHq
7T9fldeoguIq2db9G1lFdr/9k6X79tXW/R+cIMbDGHjYAQDEz8/PJ4veqqi35qYw
mSipcOQFx6V4OrNtDBy8uRdlFOV3Fl+mCsTDSD4m0fKxl29E/6253I5pDly9nmAg
0xXSGWk75+ztDNon4drIj+vif+GhoWuQPOwPtIfYDH62/ssuZUlr5uBZNRTFRAp+
YajLMy+kDfzaWmHAe6RHHiJOQXFvdyDt7gI8KwBhGu3iLXOIvwtdJOZ6HFy41APK
fzXlplZTUi2IYC1a7PAHnWxYfIYb/pVZhl2IwtWrYUv9+LCJzJKwJu+NIONYtrkm
/RO2VDRb5aTJ1zRfoXH1NSzTIqkJ0MgMWRwfBR8ysMvim/vP2jb6/THunKcllUkO
CETnRC1RwCRktQtwz3ueArisn4aqQK+XxXMtoQA0hArx4Go3aonxpaPS67/3kZpX
NdUWL6KD56YkYhXv61ig0dQQi1lWciKl7Ugd/XtOWUCnMDnLYK1xC5JgUADzIZbL
8l219X9gAEqx8AbH61ezm854O+GNhijz9fll1uJi4aBdGjaQoWNTeCrmBz1HkZOG
UtHQ/eQlaQiJrRwH2D/6VyXe3UU73hyJ/rUjhbdJ3RiImwBtEW3/fHI+/5U41ZeD
7412V0qY8YFoEIpw+GUzOye4+Le0I8Q10adyAC8FIHD6QI+liexIZT1TpOSd0Jl7
U78fxPVZRiakli8+cn7boUyfo1al7C2VnjRzsx55MiAq/R2cOq2xCnja13/oHgbp
EOhJsm6+oK7XhnPD5BOvfyfnGsvWvHX+ps22vVWI/KWOPsB62PWSZcu9LcvFtK8F
gWwyUieM9EtKDZN75BWu6b9QVWx3xmIaKwu4v2Qu9rPTPWoTG+6CiT4GbWqSVbbe
hJhFZHgBCecUZrUbOR1SMxSCB8JUo8wyTNodHsVmDtDOVn9UNEd3ZpNCQXI587vw
GzrVmIaZ85yzfjO5WgzOQYQE4EIDHpbE8mkXBojy6gmrAlSb1P1mpLbm48c0jAUt
Zv75PPSFvy5Q4li4Rc1FVYms6CXYK1UJg0G1KMR7Icf2Gp65C0QCiRMvRIxilCRy
OseG1okJTrK6v8hFWmfjSEm0iV3sk4ljvTgyPxkSBU/c/473Xe0961pX3K8svgIf
4aAD0+zrubCcbbyQ+HAtl6ec/5PSoTp18tuqxFHEELhltQ3ROxthSRPloiJ2qcv5
Sk+/8TWrhNL07oU5iemXiMlfgGcg5boNr1eTddzwp3lX5SfCFVDL/8y9SXI8DcPU
8BqHFENupEL0gBCKjL3nrtAH/wHox2PODLVn1d707R/bU1W1dozslk8cHWaa6MBV
W0a/S8YWmQ0EIHjJH+9nmr6ANXEW2TecNWG33g6bc7qcv5VmjYDJ4lzfiyxtP8El
cBVIzpbRA4n/TrURbHKDdv9ZTPp1YYDAHrzCX1EHKtLNnQrBZE/WU0gpbnuyZRUx
yWebvPrcjVLErIvx021weSOZ4I0nj1RSQg/oU5EB6fWx9Y1AA5qrV2S4RJ6341hF
NbtxbMKnAKMNA+WYydauVkrU/76KMj4UiG/H9yJO4o4IZrAr70vWah5AfHvbsNyK
8UIhZho97KLCpxL3JlES3TJd7pSTpajtVb4+bHxIi37SOtz1qkny7zIynbgGve5b
RoAMdfyLAmeabPdT9vRqVJyby5LlzTL0Q5vD3WKL2WrrItCXqGZrkRUeiNErQLgv
Q/+UCNYbixTRf5Zec1PYMugZQjlRxv9C1FFjPb/7zOZSmenlySNJZU7aStAflt+W
n+3tPeWrRww9SW0wrNMyI20MoS2Iu1wxW/KRDmyWBNND/CY0KGlmUi+VQm9c5xLL
XnSULyU0Pw/s+GfI9nqbUcYE30a6LL/XKAkfircSxjb8Z1/eCHygfRv82qSmv7p4
YWXaqA2O2aFaR5RlkAsQ9A7LKbEiRvkiQxCujMfYR8S+OYhZVWIyD4UGTLewfkPl
z+xSbn2tW8VCy2/gmUo2+k6tzEawYWoMtKZBZZghBoaubEf48SmTZtxuoX2Tmt/U
ml2NzM5BlwdYuM43f1upHvkmctBo/iQu850/Oqm3KvatqjthqxmlGGmEeYHOZ3vc
b7A1/k8kYNfoEWLtDz8Q0Bl8OWQcUbVV9z0DmhEmqNwBul5fRiAVk8HLCklF0lrn
e6d14Qmea2wo7+7A5rcAmIJvunyqLX91ibae37qf3e5x1JR632MJA4Y/nvnwOqjR
1CVw74rlywX3ObRTovV4PUb+riZlwtizHip1agjfO2YDUIwe4/ljwCbF2GouCXcW
uPCK0WwtqoB1Xc8K0U1MzqObyk2MLJfk7Q9w/vQCiuB2Qwi4M9Kl/y6IFwl4tqzf
X53O6NKJBMsj9bnJyTW5aewndXZV6kUSdWCBjefhrsMe68re8/i9rNfrQX+tQIN1
AOMPEYabHWXHQtsqJjByGzufqYul3zzjMI+1jziC7VAot7rJzA4b3gSbXltexZA6
lR9EBvAdtsN3ReaST/eTGOo8iwPMyaluCN6sQcKW2fXWRP4tLNxFSTBaHlJFcMbB
Y3IhVuWNr/t2wAh4YnaIrXM4pRjKI6ByZxkM9Nrtwo9Y4tHRHXoKlHdgql9afn86
mjpVs/1FJASEde7SgejfyYN3Z3n7V3J9H261DM/H5dqcT7bk2Kpi7pUOCP6/H/tM
96jiPNdDPAqBZV31dqipLuotZbKgmNS2lDvGzGKB7s/iLHWNLUTwHmhNHrAYAdbt
nH6o8jnmBuTVg98bOz+JFWDJaArhXPh3CiCWtgSCPLm3Bofo5Fz/DnGVPbBVFhMu
bToPl7gudImVuP7Z8b0fVn1Y5uGU/78P025zu5K7P9hE2zibr1q0ZYrc9ef2Ybb6
hbqzkIre2A/8mHb+MbP+T4dtTrV+qVA2R2G2vGPGBcWum6dg/RtY+23OXqV+/AWM
/4/14Vc8/7fjxqnyEa7D+T7lUcCUj3Re6WmiQvbx1myGWy+l62Bd5IwIzuwpS8x6
BUYZxQDNVaeeCXzbyxptBvWDnbh3czRRiXGg4vDxmmXYdl7ueqlD9S1g2TgaoomL
lYFAxFlXHbaIIpgeKsAFgWzztyDUAa8IFbMhJl3CQYeG8ro9fvnvyQzXqg3iTdPK
e6gLHge/Vz0lqbGs1UmDwsuQsiyovGelDRwM1rhL/NTEcg2kR1PaL/GTgUTnMnnp
u6rNEiJDwp6W4+towL9oM4lzhUM04ofyWo7/AKz5GXm34vDTq4nPP/F4GHhFUMGH
UkOcTDmJmP891cElk2tjw9Xd2jf+s8oqOmDGeIel+hZyikfiyAp6sf5BUp7DaRR+
mz8DxkFVBKfhP83ca1VxS1GmLPLNn6bkZ3t8tlol0nPfn2KfoXd8E0SLYHSba7t+
FSvMRvuWPClg8r38aPmOtdwyuKDVndd2xOwGnSCD6Ui7MG2GdCm7H5eBDpug/NvV
Sa4V5l0RTeerHfiCIpMsp8vDR7M57w1Tf5xCELcbELl/2wTlIu95iSW0H+M0jWX3
lasmeRYNUflxcFXO9stHZNQAD1G0pSJ48rFDg848QQRJ+4sx2WjWj/z2NTx4UWhQ
ADhph+584JDwECoimX/bCic7o/uHZKJcNn5ZRGZRklAtO5Qsr3JhnnGp0ybgghTc
jIQ97dKOtk7gpXyGEn21FxpVlGUrYq2XAYKyH/f8gkzTT7/6L679CKV8LpTtvdpM
6M6WS6nYUxAjaCCC5qPekUKowRdwtreLs3vVjvTU5eUPMCs2r1nJXKj+nMByv5/c
zZQf4qVzus4pUI2bdD2gyhfFU+0BoT3qlB1I+s9QupwKAE23/OsqEyMFz0Sj0bwz
kGNhQ07YVKZfz7za3Vc4fVzUM9vksAGI1vrRLW06LREFkxPF2hRPYdMqYrEepLT9
oc4nyvS7d4xPS4gUFWlr3t93Q8J2nMwJk5DnP1+oSb0di89ludp7haXlSGxSLCiO
9IE3/o0y+aH8MBBVvsMAz+SnO4suVWbxeSKesJyjbBkOYime4lSCp525/Z95o7OC
Di1020kHbtx6jAR1+fJwrskXNYVk9fAdzImtK5rEOl9bSM1HSvI1rIY3Gb7eLNWp
vsGDFO3eGlimXXHGrXeetnCTt61bv7d4vlh1A+floZvzMuaLgYP7pJFd9HkDl/z2
eKdAUONjFaVgmuR+hxKyqYO8fnOICdwRXKMfgPnAZ7PSbPHzdH1OsMXzRJMFoRpi
MsKkE1oe30LNW8Nl4KI4sa5YIuKpB0wW2hE8ksqTJaNTW8y2JSurhpw1hd+5636+
2vBPPmT8/12EU4nqg2DpYSCU6xtRImrE9TBoQA8jLHdh3BQXgQzWi1CeL9itmeMw
opKhIE+6oJpd3pVXxkB58Szk755KsCVgbCnZzmhu8iEgzM1v3dXn/Sb8vgY/uQKy
3eJYLtBS88ur01Fc3xgWbnbBdiEegkUesROp7J2O0eO+LWOyzFfdUobPrFw+91jf
aJM/IoPazl11HlVWzJp/24h0Ly4B/VwBqVsC4msJy88edAeiZ3slSRrI9uunZOVw
EaPGKjVNCpvCcUpiYnbDw5VT7oHljglFfPSY/cdIhPL24Kh19joX4s8KYx2nW/US
6tS5QkWKwHZYebiEDACIOorzP6zJFgd+xQPfLwkPkQAzel9q1kbriX/utYmIF/k/
4WC5ahOmcAwGTOmd3fadBYFe4McEmvPNjK9YkvFCjFEuUccoDcyDRMDa/Di1SXOj
0ePeNZ3o5jnyez/wyF0vF7CZ64Dnp6+D/vYRm5SCz3uOZIBCQ5FaNprIVZjIJ81N
RjHuyXB78/FApiMyf+j6FK9+WVjpv0JT5fSdiNvZS6cpw16xIbkcuy5vOI+OQtAZ
F8/Np1RZ2WQtSabC6lDS40sAmrlPCsPyaBYg4OzKS4wValxfBaQg0ermKqOV8Sgi
HkaFgsrU6b2KALrD6ZTZ1SyK3XqiTD1rUM+CfLDLEJ8nYc17lVUoKQgIgJBFMvI2
U2Gj8V02P9gzpW6ZM9qwzzRIxK5k8n2JxN2+62MbVCpqi492jszxUUIa6AF+4GqI
m3OnUpew5ZOB7+kfF12+LWGttAs87EiUAa4iyqBVadFWuQmaNYpvSS0KeND6oNmQ
2Dql7xaZXgckrBS3ZSD9iUBgaMLdVukQJ/evK+5P08g4k7tDiMmcjaF75hk5S0Us
Y0hK4YHskXuWHrRT8boWJTvOhh55KJ9nF+Xv/dARnjCp+U2yW2pSMJMS0rFi7i/q
bf7MirD1oYUORy9fLp88Noizv7axx9xtxb8CIpRAjCZ3/e6hG9dT+E10ItNjYWme
muHiykHqPLURK0PhWhYJNFs/hmlcxVmunIELphiDO3aFIPzKHUV5TE9O/J18pgFp
zviuEUJgp7gXn9YkD9YoHdEZk6l9YD29Tks/YiWrgFyYlyrjzT8NSiyDvd+QDnPc
V6XOCccomBdJXNUVNAnRMrYXxI0r+Z0Oab8kYaI4KJ7J+LQvv7eCSvIQNVeWJIzv
JC92WnTe3eXw+Wg0bgMpwt3LdqTxqg43B8ds9zhnqi/a0NDhlHsHISLzWWKUVYxB
lXRtZ/qndiA1bpmUb6LXJiz1cJ5PL3c+kOPl9i3I5Il+d+FLbT7UvvnRK5SfmjvX
ddX2BiKqnY2YOKDgdOYS0BRoahZEpwSeDWUJ3P0BMYdyHCvJ0p8uylm6r9MdiZ4h
wvJxm6HHQX4abU2Kr2Brtjm5YXcv+AElSwvwKzSTTWbKtoHvxaa8HpT4WZ+zy6wX
yue7gpf0qvLPBGKFw/2z/ZmAmMBFGdgBz8PXAAxY06ogPD3bDdGJhdu/IM5jg5xa
XHGw//eDCI691Um3rrl8ddhRMxZuDlWvzcJOq02ONpBgqk20lrXmygc2vlkIt8cZ
jYxaaFFEn+cToNjp8T8tllO69V+icB8vtOQA98C/Gw5HBFeUjMESdZ7kzaSbpuvV
lqeXZUqbc3hfPMWS3+IXShuETsv5CFdAa9uj3ydr/DwlSAfz5Eei7r0A9TVtkukQ
Dr9156LfX05zDk35J01GcJrUwvMrKY+/xpMEc2llTArT+YkWK6wufUSQ8umeeGUD
6mizwA55DMttSehN5GMfUPGdv/itXW6ezpnCQWoeD1gfqBB/odskSEvHokO0Zcar
QaTaWhz5jPHpPoIfLxA9FaSrNUpgvT6xDpcuNT233bueWWHnRyiwuhdrZqqjTvZc
HoGcnsI8blgV0JgzXfVecsNyPdvlMAKRUyjspkwyobYGzO9IY40fGSPtEeF29G/f
YILRFKuqCcp8FSh1lZ9MtYU60pxP7Adcc/zWx+/vT1KOGThPopqMHYVMkHp3utJ9
rM/8Xa+9p4mQAl76vId1EEf8jA7QiTDTm+g2eUJFYEukY6/tujUEcK+eSRV0GxY6
Z0QbucWgoyN2AixkNEz7rXctzqk34Rrnb/3lZc5ZawbnE3ybMDaSrF046LDo6fLt
NWD/b9BwG8sTomkpLMqdCjmlfzxcjPtmCF5ugAbc128Yb3YReytmnbm27viTvw+o
P63go/BT9hqHpZ/miM9F3d1YP4Vi92D+Qis+qSwPM8mDVwSZnmvqLEa/YgTr3t6U
6LqtEKGQbPck8nwT4zpz2xt84VVfkaWLKTjIvhnGIEVglWg5niIN+/cwozEybbHH
s6tUtr9umypeoEaWeiOBdVtjogJR7NhMW9mUM1YmKAjVKFZxbAmbQVYlRlBPmeem
sMWJE35V9LduKoiORJ1WLPgIuLrzc4UNPqUGOsQallBvnv+k7p/eq/iqTWUC4eCW
ofLjTE6Np0OwQ39wBIHvg1JRFbmXkYoR1eDA52IK7zR1d3kJD+n3QlAFu3WysR9v
T3Zh2vJ6eLIq9+fOUmbJMi4S4EVsCgygfyHBHERblrycCov0nMJjQelBtYrmaOXx
YWOcC69Thr2D4Prm+iadEPVpvw66OWxbWaRZr06tHcUJYcs57wE57ymavx8qDHg/
fdQX04XBVW+3dqDf3as1ckUmtk3VIf6gRju36rAu1wshZgdJsq8zQrL0jiEH/AwF
C0do2xWtW2wWvdtg3vy9oNljJqL8Qgrv38bOtXq+MtBpwHX8UQIaS6145Nmr31qD
BDIWT1Jm56gZfx1cwoJvzoQqyGks1o+O3Ko7d7Zo7xYgIOFV4VfWEsW4852ZuOeQ
0q0Pro5nMAXU8dVAsAJcqdP7XsIUCX5ICiLHBPkPxYgyQtn2J3Z5inq2IkrHcX5a
yRvF73AWPP8IyeL6u+ewoC5iVWJjafVxXCwBgquJK9bMDzIFKckRnXAQSmupa+G5
nCBV5HYUwjQud3DEn4XGm7uylFERGbiLxQdJ8NtAquypswUQkPxO6t+/pv8v1On8
dIvJnCf/dUyzSrbu7Jt9IQBZnHtKkSa9jguwmjpUswYH7geByfpwLYLdPqsy0zuw
QkIDOTnyjUh4XmsVZCQPkp0reGefdVYbqqRiUpI+LBBsy0XIF5hQWZSjaOyXTmok
RKWIw6yjrSpBHk7HypZ2XAsSByJ3ARVrM37C+sh2KZSrNSLm7MOoRXN2J5O3zeEi
coY2+0Qny4fMdycS76O8PMTUVlGOzsgWLPk9knw8CgPexdeVzsxXeYk2hnKPW1oa
d6oeM7vfkHJQBWyk00qLfxm6Wiv06RNY+/sa0AhsKMlx7ej+rcVV5sv87hvXMy65
0SyECJNnUUdWTY/82vL39P6DBtkNL4oiozt+eRT110Z/H15kPrzFjnwuMy3xBv7N
6X9FXv7vvf91OyeEFK9SGhey64SE7hU7u6yOX4eg2oocu///yc1Ae+Uyz9mA1zNi
YPCeuC86TPzy4lPn/QLD/S9sBdEIKjoeAryg7J7O9vPSE9k1QQA2e4Vc8Kh14X53
gmtgxejLvV1RixVb/wroP1x0T1OKF/huppu5uQGBeay1ZmVVnNnqBzzvzng/K3/g
2chYGtIjsvGhwZsgW7jwJPrfG0PI+GLqG0zVjlwx77zGFivLTngfcbDyAx8zZ2A5
F0pL5jSB+V9ok/Gm3xzQiDydrwIvGykwXowS/S8/EEeldC76OmGUV5GeyXHY2Q19
1iN6s5dXQTAw4rhmQ9LU2oIN9sY3fkBgNSEkaBtY9w8UMiDvsF90jF+yPp90oIFt
uIjGoJUL6WH6405aAeCc0Y8HjIMaiGhpf3PkJc0Cn/DcfsdDtjx1qfT0UbbAXW0n
4Neudj37JCfJRkk/3jkGD0zpcUxjFi4ZLQawdX0ajmIZSVK0AVxoNJ+2nXgNvFjM
gXnJS4WDZUo6KWA3Sfxt/XL9TdQNC2nN9pMZ9dn9fAg40fO75I19ZP+OqYl+RgWE
5wHKjzN6tpJU8gpbzFqMPSB+b75keqN+RiDgLbG3M7jrH7WFBtYMNvFIya7jDnkt
3Vv9YrmJMPkCL9ErTzGmwTULODhskh+X6PlGZAPDoF1JuDsVvFZo/JjT66jXkq3m
es/7o8auYYVB3shl840XGEDHuTmNIwXc/O/j+ucjtdBtieuon44vtZaQ/47hnDh2
iRR0TuDKaW6l/70jP2GiL5gfYMFbHx9v/uVbDg8wuD+gQ77vfpHqKX/yBMXg4doq
BmuUqrMu3T6Z8DXIRdkeLPa1VYJKLTDn86FFU7msH+0mlkLs8c9AgsVg2PbDj8r6
5bhIl1cNkZa+8Jz2iJIt9ryPRty9bbRJBMOQjlKIxE6lRn5UiJ8skh/BJ0bNZI0S
Zru8IQ1ohfclulpcH50uMnHsXSmXXPSHhxTISldluCRsUDZ+qigLqqRLRwkuYo+u
QBsE9HUj4g/tLGPnh9jpKLRRZyZugk3+coBs77jMNZ3P3fHtHoYiwKPg0b5Chu7e
wbVpaU427x8gXhrSoOzUgrj2I9R7OPkLbGXDIE8ohptMgtcdPbjY01Eunpf8b1c7
E6XV6wbHlvgJUilMeOs9pFO2mFosorl4ryzP08vleX1Qk7Nxl3QYMynh3lOn1vOf
m51bNnSluTU2qBApX3sdI0ws0y+E0y3XpBkThxpKZc2Dd8EfQkcV72qSVnw1TxQs
Ayr9qUNEOdZLYKP9Cb+SwKDyBfqAJJbM3JZ+zrP+Zpftgj9VVMyoLkX/IWXtJrJ1
RFyW7PV0op20plcZZhuq59QmO4g9SfpYCpBTTKhjVdIFaWjUSYB5i50MD9BpSI0Y
3teB4bndj93INHZojoWnT1Cf/DULNJGPiJti59xxTMudqUiiS+OEF0ID/vCTNP1v
3G3Bn0LbCunMtjopkpfKen4UQdEi0j8woV/Ozcr4i4JDQM1KFhE6JJvUEoBcBfeS
UjXIzzbJ66xDO8Mg5xfhyJvH9REqgjYigUwlkz1GdHdd8b5NwH75WfUgpbeKDJLg
qSylvBgOVUkHBNB9bbvLsQoDEJaEmOpQVMDa4fm7C2u3cgAaVaUTmwA2iyOTQMUh
u5rw2Jxhi8BUP6PV8f5mWpC7s5XeC2CZttdHe2UloMCZxYyH9tu9Qngg/a/mL1wn
oV7koB+/ZfJaKJqUTOgjiWa/zVMYw32eMYPM1Cj1Cub9ubiHBehipV4UUPuLQvsL
4LHY6QAyx9PQRWevbBenTfbljL2b62it8k/HCG3n2Y2lgiHh9E1+W07i75hq8gss
0nRpR9aCAmihuhJWOKzlkJeAHrZZrQiyOZ1TAj2O0Aptah0L1/j5Ow8RGjDjeCTv
Sr0L72pSq4abO2fcRbxAXxkj0Hy4OeR9l4TjXvJdNGVpdIFBkHvN02xKHQYM4WaB
OF2EMUZjcHimN4GmDl7MeeuvI4tmdep7J07YyIVsSryylQ2W00YRTLo0Qe1SznXh
QF9OPTRL/dzZbKmsd4yH2IFDHPnlfsPTgkNxKQ5v11ASDKDW14sP9asmDwtgW+Zv
eCDgDWXg7rvGjLweyqUguVodOvo56xhLpFfuqaF3I4Bi+lMbiNtyANioMB9pwuMt
RtRkbSuIV3FOw6z/5s+7JRyUpRtPqIin0usmJxuCRKEwb90WeY3O8mrc6Pp9Xwe+
+GhKnMK3DW0o0J7Mz43CivHVJPMjCrz8YviDGj/QW7pKDqEFH59psozVJ6dNfArX
Y1FPVZSoXsRNmZ3Vkis2Cxm6Y5JlV7gcKF1ijNZJtNL6eBbJwrrZDcfNJw2CtY47
6Yu4jyjmjhRLhmYkZYgC65LN/d7Cf0r6+qlxpEwDusEkXtvTbCVAPbpYSxBDETPO
Ly9DVwoSe+tmNoWTH1bZua3/H+kDpljWq5yB5YYv94TlyApT3v/nN3MfOfBWRa3S
yOCYd4KngJXCqToxRxLiwl2OLVnar62ngqgEF0Q5W1f9tcO8NzyXurLa/75EZ866
WgfG48zfvuX1ocHUKpKec7Wn9rdRDTi3w/cs3gQae02Rd+0+U7rRIHDpnhp2mNTc
//bg8/RwEDwt/ecO0pTNH31Ka9I39cG8h/O5PR9+RqJK5BKhKwQgv4NVXPsdI86x
wZMNB7S4L01jkTDnuOzS2RPGZZu8UVq6tDBJABIOeZKRO7yldzPnjMnRQ5bXXGmJ
B0U55K+rX0drHy+4QQQvkuvvTD7CRWlQkPqHZw4BfQ5pzmyGUaMjM1dwupY9YjiE
aluDqEgM9bn3XFObF6fjf4WxFeRQ16tQjCw3vG4+dn7zpamZkJfBlL3HVrWFysGx
oShyS2nxn7vsw/SujuDa3s6zeN1UNE7paoWpvwVFTw+TULyJEbO8XHJTrt+EoYEO
TLiD0Pto6PdujeJ85FAjHAmb6R19SaFJTRCJSihjt5gC8S9mR57qk+q17yN5Nbat
CylBYuZltqlgWKZIGhDicEVHNzSVT0pMU3GaEkH5WzWdLRwQHNRn3QUQK8E3SOFA
8PBdOZeX/45xqOBxpLGz1jnU4S5NiirYz8Jclgxriwm7sBs4NAVLitqOU+4YWksI
qqtp7AM0zbHnVXbs9Y4zzm0a3usW0/NBXRyWe+t8TIDXZ7KOi23qVyGB6rwGINKf
jlUFWkXIOAR1CkL+YTyQ3jvtpO5ANqDSWq2c0j76oPwJ232zi6kUv3qkPdHb0C1S
HwGOMYz4/7xfAQjrSKVPltR7Vzr7ikmXg7HN12nUQZc/4dGbbE1t0vLYag+KeiCm
xEhlcf3qOFlNKmxMNeRXaAglgvHJmi+f0qElKCBDWN68uImPq/zR0Q9VutjWa3h/
rGH9wDV+3XDY9bXaAiSF8WRK6kO+v2EhIWKRqAhkNBJeU2Sxm3UcJg8DUQu1A4Zy
ch7UB0IAS/XOVVnmgTD1kQdFVCtMj2BlYGvAznc9KRNOG60su5nz6GLN4NEKD6wq
6JFfVx5jFvhpW6Eg9D4ORdrnHXpldPz4h4AQer2aTPBzohYpUJCrCgmNLT0Xx+0q
2+VTDlWGLCDMLNFUqW3nCGK1iWsHnKuZS9tikeNVf6jP9jW/wlDoY8Lgr9Oh8l4E
wWDFzTWSawQ2mxVmoi2ya/jUzwZLBql2Y0tGrNEgLwulU0Hk6q5rDvqk3liDoVTg
Cqs+NWEgfK5EIZoSQZla/R+1CMHGo+mAoKQsflDaFr2nWGUZdpZFsNRpQG1OwR6w
mLWdRx9jpkHh5JXYr/Kl+YWazIyxNB6se4KYYq1MhB9VhWgmfZPDRpPvOcrC/AAD
cvVSG6fFbUgpCVBzUd3yOHl6ht0HpBTJg/bTcUy8tjhdxd4fZEGZzr4uZUBpQx/F
6/qUCve43XN7/eNWPXAKeWnNiwvKmTgru74pXiMhCMtDmqWDAh5EM7/ZUdU86jDk
mEthIQt/R4J9N10XFu/TTylbVMs2gKEiXABJzRUrTKuVIleQTp8zSn6K7OjW742S
BaYJeGTLPjmwas95iUVumWAI+CxX4O+NfTd1RGGxm62g1HqS7EK14FNv5PAXZDY/
+o0Z/HTL7TF4HNtNyat5rYEr3+tXyZApOY04wLkqemy/szCX1Dn1cRCg0OX700iM
mO/LJt9nMIPwdIkxrfyIYhevvyVblZHMo0UmtrzK6alk8TxqjSV10XpfEkV7oTQn
Rc9uPvkN/OAhEhzH2FTjSSxQDieUIHHzTVTu3onc+cP8M8c/RU+XRQbUAcnkA+CO
R/V5TBh8JVNXmtQdgJHtiF+fgd2LYqWF/1r2/+lcTsSBRYeino2LfjHKPbw3Y7OG
LFOKSJV1vzc69GasQvcXpl2BDWuifkAvAst+xm/KOBi+DgQ+xP2v2/m/98saFbD2
vn/Ml9VOe2GgU3IiNa0dyduK3mCDuE4xbp3jjAP6mSz5zQRfofWHfDMZQEL8hCC8
qViS5hMcG4YtZF22n3uRZ6UVku62dRHbvs7UhFxuMmQUnTvPT6KjSangxChlYZqt
Ja/pFhAwztmra1Vf6Bq+1wZJpzFfTBO5UsawJMLP5EkudXFWKRMbZDyXZ1WUzSXz
wzRKFCt8BnvtzT0Yor9rpntMNO6MVikfJTJzDhvnKsvtVQHsQwflgX5duqU5BqKu
ysv+6ndiQcg3ZuWveKH/dzr3NkQxH5x/9/Ees3JExUnqYPbg8XY+xsbq3XBv3PID
LqrkiVzo5NGLGXKjrIWZSBQW7kC7wnzwurDdurok7Taq/SZLHA9Yc99+2SIn/PmM
E0jwSXJNB8GbZCezo0GNN0uCW7yeaQCDkDvPX6Td02PG87ChxRTrhETbNGLFFysb
Z4viFAkZhFj8Lk0IIFRXtMLItWwaQf+1VpMxEJme649Dr5C4vTQjBA0jwDFyWJyU
mv+pmStcudoz6f7l3Xo3uvdO7lBbTGqFVkdsCgBKC53BJDQw7CgS8dXMFcrB30dp
GLFRJPefz0qpSS4v1GsuZJFgBMZgbg0ya2MNJuaagWybOgJVZte+nl4Ugyba+A1v
ldAIyc5ee6X83aqHnsTayYEJJ/iQaZK5kYWHPAKZtxsGpn8PRXeKQ+uNc1wa65Ub
RiTN1JJB9sDYjN8ehYA9PPyKojDjFl76bo9iKHcTsAGlRh+uHxTJBNOgWS5KLzue
A9SnjlWG/u2R0YqvxTe5pPhiWPfUFvx/Xl7utGhSLjtRpWyJX/AZtSPhF03H7eo8
o9eVoy9sCGwCDvy7fdEy8M0RU+hq+A3C165xhmxBr1EEjIT8QH1T0NNeNyBcql4z
RJ/QUlmcZcVWTluDFTmdOk9gRkXgLl+ABAp8hc/+Q6kmA+CO3+ub9spz/3/B/kXW
dLI3VnwtvNYv5FgYim9E44MTSPhsbXQiWvH49mOuwiVyR1qtEJCUN7cQJvACThuJ
KFzsS9D3gk6hITPkTUI3jR2hnSfynQ4iK3IKusCs+sMPhVy8hHAoa5NBhrLVascJ
sIle+vfzWFgD2H43iApki+K1lpo0ZZ4072c+NprZ66ux0wyEu9HRm4EoYef9byxu
8Z+0K2F7Yk2eMrfcUDPTX19j368onNt7QgFCq3+JGe6i//W/BF/uJyzbm6fiyKKX
UkKM4w3AC4DQt6MYbeX5Ugy7wIIlBowu4Q58YByAMAEnl0XUF36vJECP0xoZugti
M8qZ29n4QAF7vsbwhCUBmzGN0iD9fxcF4TNodyL3nAGi5lF/UkWnYWCSf7+2YjQ8
bciNbPPfS0oXk3e2fBhf8hRmV4ZoWs1GpsjHQhqq0rj5rRaWYhrhgRVS+cQEHn+t
/ptj/BPZhyQiv4o15DPUoYKTV+WF8kPafgRQVBTb+QVDR5rfOt9FV7tDJUlbRsWs
nlouxTBis+KwB0LqACHMWqERw1blsT8S73JSzaHPFMD+KJYQBa2NOiCiUm/qW29B
bso+AkrF7G9zZq46nt+OlVLFDvhnpy1jy7ZVWElVz4GCnJRegLj5wN2JMZtkG6fS
Gv/fgAlcg3SI/kKaf0Lx54tVECmOzb9SGHCmHWoymp3qMqsMNvCvzljQHzrK85YH
akBIqf+3TbApM4p4sBWF9EpOLkcqOeRZi9AqcMD9z8j4JJtUb5WuxvSoFB+6VLaz
tL7drDWZKbhU9LR3woU2fUfzZ7iAyVDqEGQODmGoei77JO894rrDZsF9Ht/0eEee
rI5VIPqFKG2UYjwcRBtarHfTVuactmEZQu9XrJnD/dHfxAQbokA5CtrwGqi51mqC
Mr0C5TVQ0MSAvplxcRRVAoMSvy3dvjHOlsji6HvB1v4zjqXZ1RBgMJ5zx1eqx02a
HLoS5+59OohHHQ3OJOR+yo56MwwrrlGm4ChshXKlZc8gK5lhhQbXhUr44vrMdynI
Q8lPmdPhpTZfN4nUeij/6n0EVpsJ8V41nzRJn+mOR1h6pjq0b5S4aStBkAb1jexl
iIcN9AOpUZDvueJA4IfRExEK48RAWYtBKWhEpBLMHq28GXIW49oDAPVqkuQgtX4s
nyBXkQBmHszO0ri5gqKnMAYHQcFRNrLHelKG0C8N7cqo1ERz5s0iczOMdnAmfoRR
mLxejIj2ddThS0wEYhGMe+RFF92SmhNYewYxKwZzKrBPiHd7Ew9JOKb/YwBDtReB
CoxyMvDOTDdlXOz66capGdKs+qrolWIKm97oJo5QmkIZqNC1dxRpC1/V7YcYyIGV
K5re1m628zS8cCye02LWLb0eLFi3oFTMkaWoH3joQleN7D+xZP2Cae7ScOHzOivX
eBiNwdgD+TMymk90qUofW6qUG3ukbyOi/ris0TiiIBWkQ+5F2S3jLzQJdJCpTwCW
0lWnJBtQ52uVFtSEbQpT0IGFKq2njQFC/3Y9DTZRLvxvQvR1OZOI4NJ9lkGsID4S
BJQW7BhBz9wcUgRHGUtiuYGqinW1cgUYUo9efu7rSinoStbCOMEN02XScb70uh5y
33EDOG8E7bFYkf8dqwVUYUjWFDdvWW7FJHrSmhlfUltlLv8MeG0+PFmJO/dJ2Iss
QU/SwloswtzrONprAptt55t0NKIRlDCdOomnak1qotaCdZ/d8Wr+G40VL+kbD/0M
RzXnuDKh7pM7cjGXfXGWDrxZCbpUgbon5KuuFf8KCR8WvwtUWHgeVT9luBOAnGJ9
vVDpYyrb2ScM/000qXS0NUPobB1NHugUvgA2Ic4nm/K6QR8+fUG2sLzT2edlS351
AkVqYL7zWBovEVqmR14I3jNkCSt9gBLtfpvrfyuq5Dd7vmubX9d5MlIcrWRYkmUL
P6o6EtP7MFW0EIkaKfNtz+O4KHkM4CMChjLh/0pW0+OLKJ+ZYopiN9ZKYYzPANPe
R2nENwtmZADkYy9ZsyCi/i625EQkqqs+Xm5cIBORrQ+xVA9BHUi7hK3UHlzKBpoV
AuA/o5LA0K/TFxvdyvblxvK1PQpOpW/gtJZDBSvCep2+0v8KVAWTQwMZ+yQMNCuy
eEo27TbEgJ75duFEKtvrFOkEhQian/j9udyK75nv4EcsyamTCV+P/YwXD0g5hvWY
m0LPQN4YFNQz15jVQs5mlohTLmlwXXslWcpzqmsp2u05UDeWMKxC7OLWc+vCOpDe
gd8AdhQa2Ezz9epX2vjEQhlCp4GmZCUCRDAH6Un0l4WD10EVl8HCgHapmmRxe6F/
cfmtMbl9zF8LFP+B7lJ9bGlHX/VsZ+f/pcJAO+CvHaQdT4oaHVbnLdGSzBv2dYz6
YxOI76ZfsK/5alsBxC3ZwWnvhX8qBxn7kOdWOcngGIqsoiH+o1uYuwzvxl2ZgYpp
VAEt+vaThBbIzebkUiSNM4p4zbe5Jy6uimV7pRH4o+ZyAge4FxMzYPm4t/QJrG89
v9c91Zp9H4rgSnf9mqadxnxK6sQa5TSoSu2pxxeA2qv8xTzX9tcDoke+rFhltuwW
lo/UsTAXiWdivwQTO3xmv7vwL9eQsbB5OYzorErLQltncYXNtfwIW/kt1RxSjUn/
FsSExAftEdL/GZg66y7a5E5oflEtf/tzTEPP1tCOX5nRJ3QhsOYuBxPWMMs0JYQO
oogdfZcERegGemWTLM/AFLivj0cVZI3mKu2aTzz2u5F3fuEnbn6KTpmbWllG+PPm
o7S+DWrhzkvo7cCSxgYF8sak15o1TOZ96YgNTPuA6Eg2HtL+7fN9KuRaJtvNNJal
MfsfU+guHUomSr58h42FnzLd6s/m8WIMCkxpFkGkvnLNdhSwAr+BG9+W5fDPRTdI
NFlTJIECPy+S5IpVM5Zf04b5bLisxfYc9He9Sxzc0IuJR9MlFW2dUMGjaqOXAB/f
a6lzaNZrxyTDi0yjeNGOfoh0EaYIff5MeCN68c5zmil1He3YbRDEz/JovOrlT8Ne
5oL88JIOHoTebSdIjT6AGdqiocXtNNUXsEsClETH+A2TbhAHYma6CG4PJjmf/twr
LxXAnOdLoPXpN+dH2Fi0X+uJHNBidnSGcioWgdwp8i2b+SPJLAygr3z2Z3INRekN
InTuwl8vSDz7RIBLxeW9E/94fxoD7V09Z5EPqaj7LZH29jckDbgw8FrBCM+9u928
1oyMOPXiD7+R98v2gWOOs76XGgjhe6UadgeRPW0b3DE0USZ+HLshXENE4NrqnvvM
eUjd7uhLWa7wVCN/wtxjLXB5gSEKZl4rE2K7Hf35WicseXH6nDfznhYAjH4onsmu
ZMmJDoRK8tAEmHEX0Bpz0mr+tK3zGX0hB9awjLgW3V71I2RSgejdKDn/SaBk6K/j
DwXCQSVG1hGnbyr3B9BrDP1NLVkyb+ybS3xCtJjKjJ9bXqHhPouYewH9JLXPLxHd
9rCBxfl8FnYJuJNehcYxkUSDdfP1A//lkEHmZW8XhiZPj9HDXSuZNB4WBEJ8ZX1j
4EOCzEcVLq1sKroPxWJ5PjZ6PBVTo6JPct8PjQAN+j2vG3bvi0pkAGDTUAnSTG9a
w/sid/QHY4O/fS1K+ZAddzeY4SaSIrhe4g5rXDH08aOJfvvmYc/LmNiNEQ8txbu6
YAHt4gJkLMYkVCMjo8HyDO+hRtDLtIDOcHBix5W0B751RX/bVOYR18GkRqCV/W+r
DYjBrgvjJbU+GFnWh+DR8G49VhrPitqLSILpy+34RCVolVlqoA3JHmehVp8zFTRT
Vrcq+wybE8buiVMpjT4Xgf7aaK9yP9cD1OLZwNLJLLsQSGWIW3YAWE2JGxhC4afR
zK8+uqgkAMMqikMtjVKT+pD5ncw566oHcKvcCzW5aegIf7gG+UIlnvgTuzQk5JA9
BXSfB6xx+UJyuTmOMTYeLUe+zPTd43OYZX5DWGEXWVgTM/c5Vbt5evkUZ8ANVctY
BIVMs9wViWJ9zcONAr6ZSzzbl80M0y/GXqkxLm/mv//yVR223wxUGbw7xxMM487v
jE9N2MaVreY+gZEGmPP+24miyn0jdPNnaiatIRj+7o92rV1IlqFMxSItSkEe9Lnf
3TPUZwHX0RQHD3a7OXJkM/rR5yn9Dnzuk59M0t34D6HijluVRTXhnpWTTVqrk8eF
LHKczxY2gXWYFLMbTsMpb/qlIETPRUEaiY41qnWP2cmjtRFbb9oYRMQR1+251oIO
VD4iHt7w3fuc9aveVSO5uKEZ6pq5LQiU2OupEYjMzKvvBTQ/likPqpz0H4Dk85sP
/F7SVckZvuBQxwl8izmjboxNyrd2lIGCQh02+WjR1Xo1D6l7bhx1uy8OIAhzk3sT
I/Xou5MKjAFNlfOtMyJMqAOy1OEecyrs5ybTZGbxcTZfcCwS8mpr+fijLdGrIPJB
hKNR9hDwHkVSAvzA6VxuMw8xOL/JKSgJqqMmoJcQ24dGTFVZNizvWNcjUmZvugf3
Uc9S6aUTEH7pqv2yyftLXSjFEEa675FMUGvGqiYkvGiIL0e41B86njV3jOUzdErF
KLe12EzPjcw6JWY6IXch7w+cRjnkTTPuu4W15VD9GUvRiKG9nYds764qKzLJjXHW
lM6MEDH9eLbS8HgojEzS80eHXk8AgqN6CFcyY8Ko3afI4rKpS1OieNIdFnlBJTBd
MNDH9w6xhktytzqewi6rSjaVkz1/UDhgMt2g+knKqfolr0PNT21w6NDR41NnsXmi
tCacRhK1soF45cn5Ipdm1bG9E3HRk5gyY+BMMnq6y8XgOkqtX5eNNVB0uqnR9Swx
b5hJXZx+R5pag9eAK8lp7s0gkEiVjsZDIyPUuxVm5x0SrWxIg7Xq0EfGzLGLfzQm
r2J41KHh4V0Caqatz+yI85a46+SJ4Va7HJr4xudyq+bJVLg2TW2dVfiXWMV+d3Ny
cbHAvVhU3wjGaE1aszCAXdPovhgq5X9BNDc4CLncXkD6tyT6vcMWrAHy73GswYey
nxvJSFZSocRP3/f9VeEc4fwdBGdwayX7da9dS+y/huUqv2wJkWlkaUbwtURLBEc9
3sDSFPz9zTasmNMKPcUdgg2n/wketjA33wqs3oOYjwhQqRcY/aZCdo5pNVKLn7FL
tkb1PppRcb8SommjuBUk6k7nkzIuaa/h6R2oFhlylBM=
`pragma protect end_protected
