// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:01:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tjTPTr0EuoDOFzzGnFx59FLkBEAGcQd9jg6ZcrExZwUVgbd7IPRqtqSrBel3M2GJ
AuSPC17M9h66TJAuKE7/yoNJCO8Yuh9z96HfLfb1Lwykpwci4/zwGlTMcRpG7Ftk
dTpEo0vk5BD/+MZiiOAsI0KlLkN5CeBIhlw6zsdLyyc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22480)
F1kw3kuVMZ0pOXOPWj52vTchcg9P7EHLNsFsEGWcm/UMtmFOGvCUfI97+62A98mp
UmpDcJ3G5DNZexRsN47mPJnNPUmoItKQM/DVom9xDE/lerOLRbGpGNa6RVXscCcQ
yWmi2YrJzz8YRJyzJjkdHGAScE0pEuMeHLtPo3psppFUjfQEUo33uDGb2wu+cBne
ehmrD1zza07fQEbrmbuW84QKtT82hmX4LkjidyGZgXTP7CCiTfwHY/BJkspwu54C
0gTyh1+AtARQ5Xar+Qo2LzxM2RWCRP2k0jpfeubcDWOE5sAgS4RRJ6TAIwG/nUaK
tWSIGEnIePLAymC06QNQQ6Ws8Ami0245IBKSOLBwx2/Vt87wzB2+pjDDUPIvpACt
JiA5RvZkiKszCw/2DdH3EXRRPzoa3valhjZLy+XmDaVEGKPbpo3fYGcKJb8HuKXj
HCIWMptiMlELgjwM45Z+Y+lbQJBc6Ft9QQtomJVhKmjjoakjZDxXFk71FAwK5nFA
Y0XuGNPahetl4Li8SjxOehj2zPiNRglGv7hTpm/ex1+Rqs7P/mvULKMbAgGFtqNo
6nt98SnfVImEy6c2KHa2kw+0B2Y1J1vcXBcWLh0w9G3H5fTrf9LGDckKWIzvOfej
StgZDoPUqo/h9NvJiEqjpuBAkvqS+HbA9GH0kVXp7vJ2fU3+Ylkw7yY/njxDM9XD
02G1qioIxZ7Atby3ZIBklTd7OjPTlmMdaPkn/fKZmaEix7FFbpUhWMyqApL+xOQl
htIs+0kqBsdmWn0jmGCyJGUW4+Jb3YBHYq0acULe14QrZEN969TMiWFLk7+7Zjjc
hkv5FST0s6s03MGGzeOr/KwbqlHTSKrmSoiCD3FFTYTrVaoj1sKp0scJzFmpck+s
oA8pTXhYsYkT9iKKYL7qN3r/uN1FmRcGlMi8j/ntL2/hAmS26bRcu4uybYvB+48w
kUehanaGk0TUfnnATuHLZqU2NEYeKCrD+RVIzuDlY7NXjEo2MBrkKEpuf7kd+tJF
KMZ/DELqZsHxtSyCYE4nwZOFTyyJ7OAfugRZLZGYnera2dF15Ah0WuGgAdzBlhdA
+f9/9nt0dGjQk3dGTTOFDbIa4uu8ybSR62hwbS1tzUlfqa6P9S8sYNtnZcq24t2k
S/aGK9hDjkEdQ1Wt+eAj+g2w8QTE2t7B05afDw/ckDI63AR7bj0JtHRz18dEGr9+
Dpn6aU+J9aief5PgLDSfmn7WnbURDRwOeJ3Gd8fYZig6AfDp6JieET0eSvhlEndx
a9l3h1HxmS/odQ7gb5qf03H19snImxoJ7iKRo6SRT1GuUJvH5TiOYFgQu4Goze7Y
xoPtmHMbBwf+APDD33Kt9KmgKMnJI/QA696wj0fJ5i6HinqWI7XpYzPpADpyHurp
YvE0k4LIlvXFH87/WgdKC48Ay7jjP1Ywawm5ivVqTTJl6E9krzXNRGrTAt8AWi9j
6ADUq3yVlwwG0dM9SnIYPbQ98nhdAIG1Vd++HAQ8nB7bY3KPdEJc4Vma/wUAo+xq
l/t/8Jh5nDteOnG3mZoosmO1+qRC4SoPlM6OLcjD5Gi3uL8lh9gXPc2U2ynGIvW9
SjOMGCzyVlTlcGWIUI59FCAvBfqbyDIS4yjpZfZgMxuSq9KTgis2RK6hncWZXomF
jN2jD1GIxfWCBIvFF1FAAJk2IOJ9ECQxQWeqNGt7mI6EDHLtVgOX7niMAQQV2qkF
q7c+/Sms5L+ltGPpxqtSNkbyBGMCLSXHXKlTSCjqt2z+T2fN6QAlhOpzdVIpQKR/
J8Awlh3MDZDOjh8nHfYH4kqXYjhL1lB6n1KdtJu+FoSmzI4vS3IKO9/3VMvW2fU/
/MKfmM5lZlcTgPWU+MxzhQmLD1q2aC7ZwAShdbpXXD3VPqtOhPNoVYHX76YUGJUi
JsD2E1zv6yIjphuQ7U8iP1xSsULtKcmubB/JYe/bwxFxwBTiECZVYpqNoA5Y9GuO
yom5BGLD6uKAtpp8JQOMiU/+QpZmAtDr0QOWE3Dz9Wonz8C1IVivbnm2xvdIluvk
bHogsrPY2+GcYAuK7lQwt9DXzmpaIjLtiWG44HWLaR4FGd1XePLMlemRJgORLyAI
qN4LLDpLFqqXZJqEKtU0Xq1L8UZXo94pVl/Zt56FXuxjof8EmAoPzcF9RG0nQMHQ
GSsiD8p+ZDC5DmrKrVYZRzc0qunLuopD8clNqrILFw/iBK610+3iG5jPF/bA0/jA
ff2P9NmO7vDqn5EGQAISfhXnrdqR2/nzGg1KZ0btSPRhYon6JTksRtE2niNkuRty
QKtD2hJM5tK78V0klSJkPlm2KMTckbR9QQdCV3IzBS51Om3JgPJ1hABfgIIUF7z1
CjbtvSbGI8LynPo81I84DEM1CYAmJJoqTLhmUyticm+7tpHeZx4Zmvo3xAwSXPJC
yYAYRSAGAgQz6A2/nEBG7rAXnCRoQhZp8ib/LpsPjikhvg+P9sfVL8h2imc9kEf6
le1VR2cidoremTfmxdrObKCrQofA7tPyLhZIUbjhmX0+6+lLrMOyxYAKBWNGeyH2
stZ5m+16Xi14wkF2qdDO68GuzYj1bs4n6o+fmvdCWLlQa4dMf+BJc8p50mEYV8mN
2YNtC6wGwX43PO9mqtV/G0KffWgPByU8mL1hTrYoGJzD4buyzZh+EBUtrz6K6lpr
EE+IRQEuNUPthBTl6jzUVUXPyvKQLKn78fT9tgA0sNHwhML1RgKtAY5kk+sWjsff
9AF3pDI7DbhI0e1E4Rtmim92PyA/AOXC4CHB5TGfRq5aGdVrpUIFpV4PmsFfhfO/
uV16bWkvStxe6JunZ2MbMS+7CrlYRN+u5mu/+Zs+s8z9ez1STWzj1U80Aro0Q47i
rbKShI2GU8ln3NkROlyuckcO0lrbuhe+9TisCW5NbpBCpqsaptZgnAUF/7lPvXI0
K5D2acdYbDagSRkTMEtMHLqv+rpKiYO+kv+NgJqMzQ7qddWZYJAU6MsI4gdGFxI5
wa0DzsNbfOKWDTOOggHAdk8PngxdTv2sx0puTLo7F4ye6waTmZ1ijbH1ktTSE9uX
895MqI5O18S2OSMdD0biZ9S6BY2UZhm1X3pc/CIfl+HNNJB2LMALUSmEqGWfIOtk
FHJuTPyaE+mzufUSMSoH165L2fdBu4W7b1rFNewpym4D6BYT5tapSxLXH1E4OlNB
W3/I6YQE4D1BtKpty5ySokVeWHKqYzk85m6v8K99VXKQrC3rzimaYxzMRrlBzQxs
kO4qNen06psDjClcLiXzxZ6I60R3VzqCdbh+O1qvXE5AcJEIYPtaTk/pQc52CmI/
3RNKAj4A5HJ3ZF8OC0MaR5kaV91shZMwKSwy/VGWxcPkl2buvNhtot5Yrm5eRQdF
K76QmRI3TmSkoIF9QTYED7XLPYYsgq+vaKsbmqcpPfJQ43Ql7tNpye+zGDXvtwaG
MjHYs99g3cJMFlbuWIU4+b7CGmK/EWYdtiqZ6S0pYn+qP5+4eotGmYJ7ngZsl2QO
xaSYqU24JOawhfEDtUDPJ6HEXrQJlB0NkSK4w8fjLpSzEuEfUh47KqD6aHJ0Jhif
K2gQbAsr/omGybMD7QA+oFgfu35J0V4a4d4Ke61Om09sqaNO+5VHTWaW1uTriCgL
fqtOYGXP+u32RXXQfNzggv8iLAc6dfPy/qVlK2T7RR6VwNLijp2Teh2oEBpGgnEJ
XYLjMv9zw6ei+l1NJFXivlfmu0bGjNkGSS/R/sml+PP61uTo0GFjByPGuKBz5mMc
C9B9p/kgafKVn0ZpFeXdADq1oAtPXpUARiB2rLehptkvWysosc9Jn+ShamiYzgKM
4N81yuxhjjgRiio5eKhZwAxmYdgVRDcjZN6GYRuVr9hpiZ4J4QQPEPdyVI6L4/Gr
NMtCgdihD2hQI8cI9VgCgaQYxR6f8xEHtUXIAHVvgWDlgsvuooMKEYi+OxS99PTB
+DvGxhgeXxzaJr6+pTFWnRhJL0kFTgcUAXbSLcCpHxHzRyCzkNGk9yA93QW7UN1P
VKH7R2tr07eBFvcNV0BjFfQtxhP7uA9KiAyWH7iBzzK8dzNLJoM1sPuqftqKWXy9
BLXqxSqxSEjjZL3dgGIVxSwMfUmTnklfg5NN1U9AdgmKvyWv8Cu+uI6FrIJGI1mN
AplW0203D51RvEmd3QMVY9iEKBGFKbkleDooCwooRmljd1Z+/JaYlecNjX2hok1P
nxhTVXIHWDNIJDkGS0ybBF3u12BPuMuis2vL8he33CGPosjoGyq8mPJD44b89HYJ
h3l/eO3i1qKz71bw2LltEQFUYgDEeIHmdyRyVk+lQVglAWd7D+Y6rv4A7a/koo6H
0ICJblqTwlAcUJ5f0BLHWWqso/mpb0qSRLiFqhNTu/ngYWU14oFHpPZsWaHCtiiK
64Ja/21yijH4njRNjAzrp9vQ4kZplyYFanTFfOUJqYo4kXO48PONTMNLY28/4Ju0
r4e8NJsZbfoAQpJfkYwaEarhKKMvdnrSr3mXboW3BT2fP8WhSu2zZrgXxP7O/qN0
CzdMQAlZNXqy/Mctnh5jSz/arcbs05KNtss5+BiWoumvQgULXBwt3PoSeqKLmYGw
VZDfwV4M+rzkp91tGNwNMDGsrAmO7+KQLubv2mpdxvGIxHUbzwq8eKjjFXAyivwr
y0kBRhIz4wF3GwMNHWJd9jQEaNRmXR7D92BW2UIUoVnYkcnKMf7oze3Z0M9L3xGU
Jl8ktYQ2Xy1673zfxFfa0gjeNmoGH4Nb5bDBmPOhSD2dc0YclR6kS582wG0bNDg0
YFyzlzS/1F0Zphew9P9Akj3EbxWoJj+LeYuhDVQTxJ0Rg7gtqL8xSbB35SXk8++M
h6TcO/uL/6xD78up8XKJ0f7RfTRISXbsMjC2HtWnSOyj+kykEDs63BPqg/7pdmxQ
eeOKrL0GxOSZGvLHlYbq94RHarcDic/3Ox2HTIJn/2C5rGBXUx6Uv7/ss8NuYTcg
jqNC/nM0GLDYaIBSnMXsIyBjACfAsBQKJcD4QsXUVmblALNiXDjwUeZirMwN5tL9
U4qcIbKSlfx+IYKjeouwRav5NLHwchvVTTkx4OyVbioc4sFnRbVCyhPVDGpFzD5e
PEaCGJnk0Jl53Tb2T5p1eHc4gnt3uW7jRW9PKNiz1j938ruJLxPmQx8Hb7VLIGXH
C4yjesamehjPitkFRjzfUfxdthZzNJ1dvZrm3e2IP0YqAlc3rvJIhMkNbyppwNnL
+G2yoYTqN1uc1zu8mU4e4u5mKHdh0yqt8lR1QgiTdRrKl4WqOMq9leKMDOZssA20
cmZq2fy7AGPKAr4+aqtDacMBnLFVpLtp6OIlDotOZg+Rg6F69jsyDWUQr2OL0F8B
gNbEUVNtCNXDfzdHgAjnfQOJwsMh1j+7WOCyVit7ypYm1bhFyft1271+TGWw/kqF
INUdr3kFKzEgbWL6ABl2GwRdpyl/p6yRywYHpeMNf3xOzJollEMxzXyRAQ8257qj
WaKsGNmAueBUHThjaHYKAUCZw5uBlabA+80+1R55Gwlx0Yr+zEFQX4IWzBlNxBlX
jYl9VyH/HeMPVXcWqJCDkV09eX3fm8zs8IZrx9Om+RsmwMWadGs8rQhlxjfzV8bI
AQrizqMnGKziZT9dHupox7R3WK/fIi9FLp7yeVXzW7K9cL9mhQJHef73wa42boz1
v7IkrVtgJrJbtiFdHVNZJbgatyGW9OWfI/uFW7zCF2n2dfBPUdZ6EWzVVEodcgPB
bGpq8k17YWri8loHXTQv1DzgHI8WUyVQxsQKa8SvYAvZKbL8ClmDYxuVmRG1s0Yh
uANJ4ncz3rMlbQzbBbDFL9dezYSBduBzui7XYU+eIleadfxuN9nZz1z4dPDQxYdA
85enddBjcniiuWRpo05yB+2+2euAq+0nDRIWP+436wAXHuE58NIPKOLd7Uv46HPp
/l2J1bIoImNiyXtegb02+gQxzxxFdPVOWj0Mlv27NcT8QWeweOUVegi4icdV6S0r
gvLfZDjFLVdq+zq/xQxGlhLFi6b8bqrySmRIYa/8BogjyazoaLdF5aqdefaB2mka
aE2G3msVObNYXpzeia5hWSeJXJkNl1HdESnl79/NiEyJkiIh8ZTchFQKQzsLyy77
pNeWOp8eDs8urgsz1GAJVQt1ywZu4LN1HZ8G8Zo0zvlsX3EhWRR9rJirWjspLAm0
gL+JgV44lqdphxLZSuTZVWpPhNjXF/fQqvuqFnH9PIaSgJ44wGkJxCCGQdfiVdPJ
vm6J708/rW8fAbMQVardgJ88AUpXRqDnJi6V2A9sYnKNBAREHgeV6TAxDtzgW94S
WCxwiWEOA9jZ3IKB5naid40azidoQ9kS6BOagBXaCQcjE7YH1NdAYZQwx56soGth
Z+L6GInxJ+99fYOypj5oN7mbhaMS6yVaEY6DZ67goVBHXJe60M3juXDoPGrZhFMr
/I9/Wve8P2RwmlddumdC5PpqBr7cPRs1AUOEOQy1yyA75Ddxtgcs1h/1jRifv5lp
r+Cx3XEmBHm3EwpCaII9CurTJaEYdiP41kZgTN3O9AXcCwhOevMDgbzsM+FBOz6k
8BOlSSrXPZPJ3VdoV4faP0eIb5A40KA54n5Fvr83w8HmK02DTNNdgkCK+7YTNsmQ
57LQ8F7e358+EY74OzCz2FBa2hw8TAjgLDqQx4I0BxgkLXGo95uGvonTu4s/+v/6
gfsgw4SoIBFE3BAz2LUJ0puzmGzAEhg22FcIwXwTar/vUbgN1moujuA4QXy3wjNl
/BUyTWVtag0rIcL4DMH+HWoDmOOuBJEEB513539/0LTIIFZuSeTT4MxDCeAni0fg
JumbJca2LIS2+8QycpeiF/ZSoJ4Af7UkgwV/2+ojqlqrTf5yO2PKW7nCAK9vK0Tr
D1S4miOz6kzFXPpArhvY2VSTRn213heKkmtubhS1q9nvXRIvq35iISL325BBLM0b
hSQT6lz7G4zn3cf/dM+Xxvd4cqkbAjiSgGfA5E6Ib+IHcPBQaH3Ivrp5zyV5UnLL
6M2gSjRJd9NVTyfjGcBHRMfKHnyn48nNMxc5oc5lWo2KPBmZRkXwe1xj6TKpQKBW
XIZ0ZWwj7i2qsszeWOvfm5S+1BMZGYg7zvfmjYRh9c5A6ZuPLjqunc5FAhSs7wWQ
yeAPGRD1mvhiWJlVt6EPdr5YNUueJ2c31EJBs4A9xcvZ/qizwhkXZkFkEMHJoVTd
5buHflyMngAa6Tnhj8+SZiXjg8TGmZgMVvKD8oKWF1WYBn3RxXJNI6d/W9O1k0C1
3T3N5cbAkLCljG1QW8kVsFzozI9gMtam0XUCBL/CR6NjDHQYGG7zJwNj1O9JSfMq
xD45L46PYu54P8vif8mf13SX6fvLM4ba234xGzATTiR2vZ9RV2W6R62BXyu+rkUT
zjdHi+ol2mim9/9DLeEus/pVUDBYF3N6VgAY6ou6dC5WLuuMBpQ6dmpc6ZEejePy
f4sDCLnIQcaCaMlj0ib2pq0Zt3apeKmcwJTPmmot408KJexotwlgZEv8ZW7sv5AI
c5jDif1278wDmNHIZ9VGYRV717O/CBsALW5+/7utxYX9WEONWsjCo11bJ/sR0uqV
aeMNq7LCieDTzaQ5jBRbNHKoTf93czP35IMGV1iDTUY6L3YKK8DguWoGEYv3eMFv
7zCnp+wzCyMtAh1LvIt2c+2mNtUeT6WUMJ78Ps/jTGSl7swCv2YbGv2bPSaje29A
vFlRC52kNXAhIc0c9kg4MpNiun/lwPK+0VbXcicbZK66HhBBil57D5SaQEc7sqWp
y6MYrf5sQHhO/8E5J7pWniPstwKv2qrLSuEsYY9zQhTvUdJG4SvWmfJQirttFx9P
JYw5lQFfK7dcpSKQAiYF3cwQHTlfHbqVlO09cxUIqOggb8nanMIr3iw1lU6+O/8d
tE0tfBUMIypnRelkklFvwjwy2XV9bFD7CKTXYXV3SPbpYLl3/5JUisVHqmd/3H2F
yVGX5qTx3MgwVWLnLw/bcD7jm3MYWH/J9wB70dWIdZY69/SafiMIRvAi4M88ILWe
EXYeT1GYGrAgU0rdg8d861ptiESe3pp6COJxCpJyfhDoGL45PqRpvFY9jn5hvc8X
vdqEQdBf1HNALjdzVEygPUyPPJVxwvSGSzwX/DNwfOt0fEFH4197xwwcgck+e7dL
fJdQKPiBPF6HbEYPaiEcB31KwD52zW0Cqc5FA9+gttxdvhSwZL1cvH2XEO4n1nn3
hMlh2kUs2sxt/V+TRQrdeaGY/YBsrKv3JuIRiadP2+Wa+BlXR/Bjxy0+JFYAyIdE
Rh/iOLfI6h5WSodTcf2nnhIKyJfxiO0W50IbBpcTllk131uQ6xTB3dCp/0eCqpFw
dXDP0ibMVu0maqC2XRtbUFHlw66OQY6Y2rBarDPILlIxnjxhaN+ejxD4hngbbvMi
H6Un/kpkpqk1tufM4n9L48sIR9G2MSUCDOiS/CBhEYdJXXpl7x40mnVxpeYxSMcu
OSsPFvZTc3QL1wid0UsNKW7o/W7h6T/mII7aT8Gb//1Ps6TCeyFQ/gvdD4UonChg
WFYH7dzPgnNac2WvMpfQHmPyifHJP/nVv/GrXFtXw9LkyugY9roQsguRLcdpoA7+
c5rY++cB7UbiFYnROxev6QVsV6JSPZ14bP8SBCTFRvGbZE4xbLWj/YIexAk3jQN7
g9SSOpqNvcQ1v+aLBIXRyxxYhDxsGArv7e13sF38YmCnbEu7JQmKsJHAQU/T0ZYJ
hTdS3boiKdEofE62g3DJZ7VV6+k0lR+bjc+xAJl43gdBZrvGJsyETEG7cptg0vI2
mkS7y3h3AvxlV5fG5NPx3tBsqYJ9VilIZMrCvodxh/t3lzSRWt1wbgzcie/mSg/B
Er39RZBNqmdzRsmNI4FDSlTdbOXZRC50Ff6WPolp9wKTj8CkMaeSAVGflrsa9ldT
pi+ojxshR49hpSLwsncIrOufdx9NsbJbvVAesbF/sxnHGYHw5XVzm0diXRrm3fo2
bzIIbWPKM/y/qhbVja8BHItYFqNi6oKXolTtj4m29fUNeINB7Y+ixXzk47y2QMcy
GBDsXE0c5cvOmDZkAWwBppGbo35mx8hCCBEPLgm0RS22r074h5qZUL5vCkuJjUIR
UEnKJ5d9r9E1RyZrCBWnwIztpfaSkNywtSJnAWzrmtx4vEMNjfL0QL5rhzhZXz9W
YmYe4P7DIwoEtMMtPhdlbe2dIdXjA4+QERtdpfSvBEKQQGUgxGF8nW+5yTxGY9n0
WD885RvH7cDu9GWcsvmVwSktWRd2Zpg0shlECeI1YnIH2/LSsqFv7ZGnaWmoYKH6
Ucq3fCx+6EqHyUEYL40wCJvVkgs/ba3bfhoBpPh/UADBTcj3yLD6isoxp4buC0Mc
spEdB5ega6DlopoMRE0FT2SBT3XOhi0RIScB0R3lCt4Y3nPfciMGLfb6dKZu23Ng
aVzI2MOkE/lqr4d2CKs12XWokpc99iU8Mo5yP4uHHuAx+Fmw2KIqTg3fd9EprouP
ILQqoRldlbmvOMSpeQQGt9XxPv5Ogpu1qc8GYI0iY0pZ/DTCwtYZcGZKpqTwK309
HqSf+GHB6//qrCi1fNK98kxRNDPoyNxY4lJ3LA5HkALMH+ZFuIHyymHgjhqIS3dJ
RpM02hVoa6PnjXJ/depOidWoSn/TxPXT70T9KU0RnaagtSIrRpATq4de5B58qlP+
dSSHOgAtw0z9S298SfxhxRT1oYjcd7TLN4AH3CTizN0gf7kmqWcl4vLC2brGmury
YAmRY6icyOqOIKAwv7EsjMzCMBf5Sffzdk0U0eJXwcrQpRdK71RHIQD9ZzcogFab
AQTMeu2dNtHXvZNVBPk+tDYNitobHXZNvEZ/muMfs4ReSYplkUEdvFsRHuXbWg0I
EthxBsyk9UqN9XceUs4plhrJ0aA1FrFfifKaITX56YaV4WK7paeO+DQRX4XQ1N3R
zdz6d5XJ16tgLOsWwagIxJ1UUPVxxWkfzuK+Js2jnq88kzs/iN3XdyRPWR2e9JVr
XRx90Ci4hn0CKYkUHWGrS9O9whVK5d7prWBEhzrjMoOx55jTgmCAiSYtN3SEQuCH
o1Rq8h9ESMYQpLLwnQEvlK2ye1fYmcYhfuT9m9vNphf4wL9O/mTC3Jh6ZpC12S/q
KSM3TMInd48o6slcvlAM/l1Pge466nWWuEjSmPP8FaMMDq2SEliBXSGCdjr4SGEu
6Vmt3yAIpqsz1ZG3YNTPGb+Bk4jabzKs1uqE1/Hh5iF1MCXJDDZcB/8WVH0Jo49h
AA/4ZgC/0z/m6Tu62gjLO5uPWlyoPZxAQnuzjOXf1hbGsTEUow7sThZcon4qEzS3
NDDBnLp1r04WIe4ySB10ogLJej6Rb1BaYyqQ+CSe4PXbcdjT8U46JNCMVJ41uoGx
d6Vs6KWmt0xr19CC4AGXPCrTTcBWXJnP7bTmNEfS6VfHNN1EMG27xssuHJEafJ41
80dkzhloDJDsBxJ+GWHzIy71GpygPjc8pFvsISGCD5gyQnceDiXyuVSnw4uZRztl
lw2QbSWRWxgGQQ6mfoFclL80GAQZq4wxGcUkXFNIWF6bHBWVdpSAPNJUN0XPcNcb
A+8a0HSTUpHQqpadrZmBappq+TChKAWfIC41acVEZqtFx2AUUz0wu582xALPmB3F
iu9hXyEYgNZMlYfpWct+qCOUZ1zkkVM/z71Qu1HXuchWFKsgrYXBfCSpSTSpLI1H
WxOANDBDAhhsenaOBZBbmwjwNED1OoMoT1rEfB7aehtoQR3dPVau1djD7EVbI5RQ
6Oz7vyr3QGEC0dv8PyXCremOfXICDGGYidIatvfwzvnYUhICBfFcpstnezKXxawm
F4HvxXHo9zXZLMkXf+VqTpZCX5pzv116qjq18JkiU3BFiii1LDBrNz//GEpL6Hc9
NtidLohVAKJ3iCCK9MogYZW+Iboo0Wgo/zj72fuL18GZQajvKrqy70bkultVyvz5
EAX7vWYuTLcQOg4EwPTBiCGuGdOnrCS7+HBn3mXF8PjiaA6GhwpsB+OHyFCaG3rD
UktHyqep/EvNWDQ78lokLtoE7h5AgdZyjFlNp+yCkehi2r+5YjeTfKdGLklwk4SR
25RBdOUKF75pKEHDV+51WFKvx0OcwLk+ys4j9/J0JsQmC4zj8gsOEZzJ5zoqmwLO
AVb4m0Y86Rt2blGJHYkKC3xbCAsTUM1ezLKpPR3sln3x94RvSV8/7Mh8SNfXXzFs
GGTWz311+QPb2wlx7kcoTWYukBb5O++Xa3vqsdyklcnj+kRtIxY6R8BPrZpx2iNP
WJqI/oBkkV8BxXLee5PpGF616zM8+iCeLG8q9pe/sXbPGqAyR2xbJeIVs++42Byb
hsgk9yxyz4Wx1Ye/JmxIwyKSA36LFu4JPyAJodU1QjQGVOdF7u1nFQ1GAGiOAZ9R
N9D5sY7nGY1afEkTh3BEzui4nT6dKKV1w6EFX1USfnu9AA5SpwPa1UWvh2/vM7WC
692u9lBHkZrKjkuzSbjUKDPIVL/d9ojPfzLSFVO4jZ/L8TXxUe8UEQckE8j1lD/8
i8LX9WiA0RGh3px7c3dNC56uA5v39dnxsvyjFx7FlW7K1KkKxmO1cvMlKHIH450Z
qjo7qJc2brF/JcLVCDPY4W/9bpopWvouzmPybzQZEPBITrzEAMQPPI4X6aQqfY+s
7/QfeNG/LyEUEVxav8WqDVULLAcDGNVnLCpVBqhiRIpV9LjvFImZEN3+ZOLvETU6
Tq3qWs3NFtCspJDbpHvjgzNUX7tH96Qand61l1YPktRtp1dfFhi7JOz6TrW/aym2
v531MQT8euODYkrs12fD0lyHVxkrpcaP5iR1LumJouMavakuvjtHaa351VgX0Hwv
Hf1cAaHSw8h0vmtfAvGVlijO2KLn+12nG3c8nkWX2vYsKBzf2f4eHAbV1udv2JJX
ptkFNtc6de+J80STJn0xC8tzwbLFr3n9mobunOO8lrtktiLOrR/ippio9pC1ATep
oQWFBATLCXyV4quzXdIoJasfcBaRXQ5O+/UQbYk/X67TmCzj2Czua4gXlxa1UoQU
mtlsF0yLYLEqqDq1kf5vC3OaMjFlDACOILCpKlbCO9Rb/7o6esn/3yIOzvo8CRTf
62v6vWx8CnDuj9SjhnqKZed8S2+gJEbc7y8K49yeOkKrtPk2HXXywhjuD5AQPhgg
P5Q+OQAAE/kCrwoe8mz5ccoUFWEzj6ZxvDhqMgmLcqsCIGTZa/R3w8Gcxcnhiwlx
SR+Wpzk7lyqT4EehoN815jSOY5WF2EZPD0nUnt+6Bi0t2l6cBTjMVcKZGGsJMkeF
aJ0H181d1RVuCLXPUfuUnAgWXWM9kGt1Ho0FTwrX83tRmVSP1HT9gkDbfsmlLjPN
HhaVPcIEvZP99CroqmE1w4ep3GJ69/VzfkhFW7ifHRip4kUsUBbrAsXUM1Q6+/dE
0pD9MdnREkLzUERzYcNPs9/1ZErlWNHOwabtADPOt9d7T/QQrcOb5B/pDuPTliTE
iOHcO9Ig4+MBGohmzMBTRPd4kD1FbSYeeQZh2tPoLN9uFmfFhVQsvfUZNRSnD9Q0
G64NJHIFnOv4UKg+1sinstKpFMnrdeEaPeSD4MHNJEC4FeZ3E6ooZxdY5fSTLGuB
VmEDqKDA8bZTU7OIMYAssJyOGD6+04GEZeAPcSOErhw9zzQJvuoW5xAsuQKJIyaj
CMbsExrlFHl8QTON06n49jcZYswqk7z4m5Yl7lvMH/INQjNxOaPJkZUoVzmh6xtd
4rYwUUFIa5MwDAHZG1kTPrlLIgVznIvOIkroXCpYOvcWycL2AlSkg7jZ79FhCV22
LQLbZG4arsnM46ikiIPaqrPLXmPbeWq+hxsqvt+NBs7aEFKMpng01+fJpej1vrdz
clk2uC5I9tBAJpAuQbvANLr0q3scW4HuV1xlHN6MKrwX/R/MXI1I6yl9q6h99ZtS
wLRxxzkjqEpNzPo9ncoYz9YMAzFyhcO9Yf8pzB2WXsWSqyi5+PP0Qz1MkT98D7Yy
8h3Vf4aJOjXihvwCawDYWAL0GIloEhcQ9a7g6NjWojNgn+f7aNZeL3NSc2n/slzv
Cg1siKlWH0mTzyc+XF80wq3vsVQGghS/dx3ZzjAYWuXLdYEgyYqFqadZokw5ji98
H17boc+yAsEbzysepEQR9l/O3JNXh7BTVhx20PfWsCZD/w7+5mNwAkXswG50OcHW
gpuapJUNiq35KKe/WJcl1NDpT84ricaxV4ip61VVTK2UYxuL0TifxPajSVdf68na
5sFKbWARIwVQcSmozubTgjuXm+YnKqV06fG/aCAvywsub2ytNX0rcSVGO/4xumOw
VVHWYv5v7mGqnnrKRUQVsJH/mGjDyam5N90clwV1VqdKBMon5Oq6rXTY1DTF4WhD
3DM7LRzU4W9JHmpFjhyjEsryplW45wvHKfB67nWmWoONBNGraJFPBxLPnEiKCt0Q
7rMSnY7mcqo0SdY58NYTb/fhrDfnYe32oVb7wASySud2PaEltd77qoLZZYVRdKZ8
Isch2XuMnAsRvWKDjsvHOmurE0YIxFRr1qtodvNwpkaGV48cd0wx0b1l3A0btnUo
JXTafRQj/4qUoslQw7f+p4HQ6weHl97+IgNUkN4nwm5QZuVYQY4peFACNjF0B+F2
+c1wzP0vNirdFxUJZIRNtT1wZe4U5Z7I5wp/PAjYutFpmlfnL3WoV3ZHgZ4y++m+
v6+7kaSiJXen7jd8CczfqNJbAS8th0uGEvafvt3Aq6Kk/9KaB6WTgsSrjF/bmtIT
2D4CAv9aIzLaRcapMzeemu6NLZkiHnj9iJoQDnZg5DajVnZtC+N5NiQjPBhzqAE2
u9ThgBcMzkaNSrgR3JTrKGLVWRhtUMKJpEFOgDKlbip4MkcHdAHWQ9cETMqNLQc2
HBCkbFsDmpH4Q5heZt7uWptUvzDaxCnraIDGWnuzzivMdZrqTegOIVq+qgLlVcgH
/ykVyKj9yOSbGg7mmt/4JjS5776QngotyhLcr3RREBo1vtYzS5a57wdGD+8UT0pP
EDi7E9kpBPgGbBhqM14no6M8tAChGHNkNfGAlRY1KBZ3Z+BuQvlmEB2Z1NRuwk4W
itpuF+MZMOTSekxK68WWbxnjxxgU2KHnYTaio/v0h63+dY5e3VhzibMCIpv9fvIi
eSiUvVaP+k/Yp8/bYSMuvsr96JX5PjxDaxfvMlA719rUka/agKIKQ68egr6fypYr
B3tcsyH/FAILyrbfcyUEi8m21pM9lRh0Mt+/Z5GRu7o8TACB5JYb9cUyz2pfUyYz
fm1xC9w9Cw6f1pXMwkasLEpN0jrLWRJQ4iPRdS9Or4CLzvq/LmMhY1gbbm79a+Eh
QTfpohxGdrkKaJsAatTlaPGNsb4VARQmn1pwZj9GzcMawlA2fi4vR5KA/qxRJkaR
Xm3qyzRX+1Y6UqNw6xLWNRcwV7L04HPq+/wP0agkBs0uYYYaZJ5sqNUoaINuHx4R
2ZnCaeipa4zeOG62cmtG8kmNRfLaYvQtBitpNOa4L/ySaFbFFB8CADxVba9KCtQC
pgaKTa4Jwr9wHIie85fkwV45Obf+Nhh7MED5UBqlfD32kdHM+Rmpc8nF4wj/lOVE
QY5ySnoUMond7AQQnEsQWRL6mt9aBN+pC16ddZQEqhoiZZzpREY1rIRs0NkxUR6O
W5lBlYjVt7HUl0qGMwqs6X0XCzKiAYSqg48ij/ry93/8Yl3AuqiVasnQ7PS2UFZ/
lidMtQwg55Z0Uvl64Vp+6bOCQxmTo1YkoYt2Ufh+co8endNTeKUOFKm4l63H9ZKl
JnmjcfclI1soPUyd0+zkJAKSMZvgEhx/KxV+Ephy/1FskOoeuNc/IXEsIcF8DZEL
IkKikVPAijnDFdJAfFYRtNrM1mr65Qrsr6GrCn3w9ilGDzF6BQWN2aNeUKpDiCzK
m2TNGMqJa71fvqAbjkiEBbtHHDzXE+F2S6svkwDM4ChWw+Aa4imCxatQcqht8EH4
pESTymBl5zrB+MMx3w0KQgJITWhtdB9Gp++xYsFI4dLXSOCeSYkhhGVis9I2um7l
ZpZri5nKtk2lvbOoAQ6qN79r/qFcJC/t+vdvyyiw6ocvfxlXtotdgVxZHirToFex
XMshWiObQhDtIaejOO3bVyXvJNX+DUMEY1xYsx9Ogp498ikaoRpUeUOzIQNj1+ZO
JINFa9HHt2l/0PTemWH3KiNz8uHzEkgqZ4dFFUTZdb/oz70bmAUdvEjIn665H/6h
hXCwLjWpWSBOrSVk/DynzrEybKgZpF6RPxnV3xKb8cViYUZMd+AkW4xZz6JaW/Bs
+cy2eb4q8hAvLA6DdkgsAVyvlu//VG/u6thiwqkf6VuQ55FK3CG50MvpfRoUx7IG
68o1C8RXns7FIPldMDM3lG9utb1f5YLjEfkOxd+Ymr0XvRraTTPpNsTHzuI8hIKC
oW5MvMtaDlZV8CBTIus2lHJ23kQsVCHzOg4DDjSmOA5HuCiqRatMjN1u6kyu6KnP
Iib4Kd7LNorzBb9seL6cGCsun2ZRKnpFP7soxQltYxciAZljwL3i6kirzv1jsixE
RzUrb9ndVmlyySkgPceJ5p9bNQ1+3x3YMUZn2i+BK8HJHhUEs7f13wCJgu1Launy
A/+dECzCoaEudN3OG6l+I0tmQXWNRhzMdjF/bibPJGAWS0uii/Mk/ndWiPe/VwkG
uBH1n/eLjv40jdiG+xh8KoXXdDosdNsWI1XLaj1g2YXy6hO7lhNdkiWogHnA+Z//
QskljVMcCHnEyjH6oqugIjYnd4MXSUIDRICHfhX7bVp4TFqfEnNjApTtDzp9mlJA
lyA/51/ePNeHptkRLVNvtXAcS4MBcQhS1PZRDOl2z9YJzSa2myFvxfutliCSgIrS
cxQv7PfF4TidjPJxiZZGHsrybXXYgL/3DHgVKYE8T/10B3ax8av6IOQSKK0m7RwM
owPjU2wjEvVhuIjTQFn30ONwhDScTy/EuNkIfTOzHMlA113OEz4+KBO8qcGoNaS+
l2JxVUKqoa3w72Krto/y+Q68JJHGY8s6uK2FVJ3A50mKWh2sFe5znBZaSRynzaLi
YX1fEkRYei1IrLXb9/1NIX89qOtzVEzMIN0U29JSc9idp28gxNvnsqVRr1V9znPV
9TQMYQ7uP5S+jbCjfPPsd1XB6T89dcX05uiVrceVqUha0TrUbP6NlOhdrImt1mw0
QmeaZJfeRqd2iI+e12FtXTSCDK/3H5qVZLhQfu+DVFJRD66vNwJPy2rCj0VEMacm
z9MVZ//Lw7cMwZPGmgygi6R+EQ74qcHmJlYevFUF+x/90al+4hyYUJ1BvX8tJSAr
q0ZzAGioNJ41aEeaDZBRv00ryTaatNCKNvPmABLa9CAgR6algAaeB1jX9yhdAkGN
Wboie5PcVP0u5kLnE5LYqA3EE8TkMzB3BdBWfAG5YC1KQkOPZPt4RiCik0YpYmdi
C7LYH5/0ng4FGjaKpsRZHbbYArLwweU5uda6Ty6TNfn/OtBb9CLHcV+CWU1OXNmn
NLeeCnhb6aZO21BBVa3zTR9jcTQUdr5h5wXxQSi2MverZ+z9tzzSATxIC+NCZC1A
Xkk0fVuI9/QqgYJ4HQQ9xRZzFjjDtseRTvyp88uo7uRyJrRsT/z+OfOxq9APlSam
vz5r21f0VsgtgUvJdpamodOqTsRQSISwzsW43icZu9Jof3ij9ZvP7qIRdu5iF0bL
DO/c6NZo3/r8j40IPnwuhWtJxgMWoOBuGibIC7SP8a7wC3b2Wb72mv1OJ99UKd5M
oFqNMKgt2qb2CV4c2vUdnrof099IYoCCsHIBbtBIesMtgWe1RMjvzX0JWCprtYx8
dK9Iy9swgf2o93PMDehROmTKeWrNqs2vQiq1uI4Gdgg0/nabRmpr6K059bLoaioF
TAs6pgbBjX63lpv1mx2A4QA/gKaGmcUtjfFeyvtuU2UiChn1OD6WNPR27aeEwnzT
CW8m45tlvEf3riHb2BQkxHHBoviQGVpv/40e+h15hbOfNYDkAzSX1iHc1JVfqxNh
lnn8YlknfeeLlLHDVz2QzvGjXd6hqG260oc7oDK3tJshnMrTipkMQFCF4dzz29Q5
qsraZKV6EHCS6HsnXKOjOnmqLQmA06uu8GzZ4D/9G80LCRRz+zhWtWTrIKWcbJ//
JQSQSQi831hSnIcldFR8A+aMZPd+Q4i9RBbQDlrPMcIi/ngIqHmB1nPsRQrNjqXT
r0iIj+v68ulXP9HzwDvZ8SH9Z38y06c9rSuzYkJvOxmeZP/7RKjpUz2jyynHdwDI
Egtbhv5bNxwl4RjFDuXoF9mUEDkBjXA30hXyDeLSS+jh6wjMg7AdzsWFe4mv5ZzJ
gJhxQAGdFV39a8e0s7PEESqw679mWbJxH9e2aDhN0f9YGBm1Bg/++G4Z8mqHqbhe
cmcTO+t6STwUkV22ufNF1DQsZ1EcPFJoXBhMHirv1K3yNRo2qSKDiCWLXZdW+/MK
oGvUZqOLvMA+NyEEqkbmqDeLhB5Wn7sQAwGATo7gNJFDXl9OrcyaTCR9GP0Nc2MX
jdzv4dUiTmnPWwXls1oFMxIM+f6WKsfRcKtbEWPu46OudCrP9sOpyjd2WiDDB5yE
xpN+EPq8/z/EbHQKSWicNFe57y3jXlc4z33A0Sw8QwdA+IV05kLsgXyunyndAW4T
tiwLYpr6JRYF6sYHef9QGW6XFw53Ulr5JQTqrsYfv0ONKfu9KIH0WeF+PiyEwWwk
s2uTByGqaFbEKD59kzwKCIJ+HdyZgKsMpgXZgDT0jYWVDW6Dj3dGe1u8Vh4cUny7
y3Sn8TAJ2ffeIspu7VjSUnvs7/TvFIyH9IirBUuay+S9NBdnOQpfd7163vbhCv41
WhUJ179TcDyNUQKcLz2h4V84fS55B3DzciFGhj3VWWO062sPvGZ6y2UFxvY0Kg5u
HxI9kRBZ66jU5NUS25iAjugXsDjOYMDx1Xv6RRwATy27e0e4q3RsZdOdggM4yL2H
qVU0npWUYRt+AHEzJmOzIZAZhx3ZJv94nyy+q58tAxMeXsD03ZljbWnRRK+L7edR
8bKXPJGNCBxy2/wrYIDBbhFLSy5ZQE7O9/YsXXftO58Gb1qyVAQg1zIdqI3ua0NO
BFELNdxwl5JFvWVvYa7IGH1G+NwuKAta+eVr6PfmpyPGqYF3QmcxjIA2i9flXyVG
hyqNJ1QmOm7+68DkVrZMJAtp3NGAymvzMdJRbInyzpIbqraYSGlHdgDf42DNMMX8
/eooDDgiz48nvWi7LanoUfpa6SikYcyj4dtngQ/6GrTi8IxWg7tBo+Xqn5TsTlWx
7TYDvTkXGsNPe371yHeUxv1h/7sDkpQVUIwVD7rHiXFQ05h9rYWR99GrW8aMjuow
ovTsEjOh6VJ/zo11gQYqaHp4ZccJPSIFL05j+ALAqYcwRrYf2lHL46+n90wb5oat
oGk2OqZkmUE79/uCT/s6bZ+MiitoS15L/4l1unj9pYGQzeVNigsnxu5vjMEX1Feq
iy2YBCRC+Uqnj0V5wKdqlM7rMYhCZ3iIqvUZ0FKGNRnM9NPo56Zd6SbVPiI4s3Vg
rXeDwZQUw8ZE96Ikb8XNcIbi0qXCKrrJh/zZ1mvlI9ithZjtCJCXtaQr3tgXePJF
d/qmgyZv9C9OlLJ8CQXgfx9+UwqR0VvETjLk/C1Kce9hISiOHpaFl04zq4N/Eytb
VWbhZ4ALVu2PrmsEI7QZ3D82qU9BEjmHhGbW1TwANEGF85CbC7XLEA43tTuATc8+
8NG9J5QYBjcYVt7D5os3GMuBg3iN/IGaNYYcmHLPrff2f02B01Ezm/0tWPsjGXCU
DUWBYdIV5Av61rF7Vn+O3PsyEGXN9uzbtpucSPlfeCoUB3Bj/5MVVDYqaJkwFyzG
1aN6CF8Z6oAF/xsRA4bN1kqgYZ48wxxAlKHD+qTYw2ive+JQx+xEZXPMNeJ0PuaI
awoAya7ADDOH6HsCbA6wCsybiwlHB634XI4xp2Gtb7ArnniCeRaJ3xk3QPdJLirE
B6Gp+RbhJ9/af1dYLZNfdX4kWOsg3hYSTQX+Ms3JJ5XiIAYONY+M9Pr6qCvO4rBe
nEVVgggirGzdWWgKxvpjdx+OrdYOXCWgubG6Z2EkP3vpbBCNIZU/GArszIxwfS+E
gL1XXSytHmHaKJ18ThwpxlEyJKMuTRbgFJmgUkGNPUh7JrUhaJ23I/PxjukQ5/jh
7LoFqj2AAPuwdMILU7aEkqi8Canafmsi1yqEr3923D3D3Z/PUqwM9AG+OZHWmJz0
0VTV3wx8bA0FgiLWSvyAZARWqp7iT3TNGnb9Sm+PNRC+n7GdE4T23F6XZeyvDxfV
D0i1Gz36WmGGYk8RfNpLj+fTO2g34iZF9ZIMuQjgber7VEtpdqCJB6x6UcQGjjXk
5ox8d8hcdi5fOYLZt48zu/43Fnygj/zp6RVQxnQdLyAI2LIBY4oMbKOA2C9jbnTM
IeXbU2MI3cYyUV/pklaoEM/MWwQD9/58Jb6l3H/V8RLNilheT2ntDLHJ7zZ6jE19
E8iFUFBBIpKf/szCRpOm+Tf4yS5Zj+Rgb4GU+55ymuUDmyAKJwWJoUgMLb3yB1bJ
vEYxIdyt9ZFLjWIV31wxZxM62al0r6rZCYa7MN2mH/Wbeh2g9CvaTxvm76eUrfJY
pgd6i6NXCKv9WlWSrw0KoelndDe0gnOUkNYj7EGh42aGbv4k8KES2PgOR+YZNIX6
9wN9S47dusgICg9RpTYPe4+3EuRxcK0vjqhetccMoEckuruK6DbENOnAPq+yhNi2
8XqQzREykFDvuPkDYQrb3XOhpmU6ugW/aZfARNjownuNrlr7UDhVpiEqr7o+xkQ6
ivyqcoBgnG/+lhxg9hDgyxIwytBtADL5iVQGIPndw7S8U6hlSJ/Y1unhgmKJvgix
HveuilbtXbFMZVbDRR+RwrUVzOOzyCNrTTF5yDEM1FfJy2KmHnS17Je39A3+Mo8X
uW8g2qjt88cvZFSOvUHAIELbJ4+UBZuY6J5so82El56tynSx7ueE5NiaEsRHzc/K
LfkAmPPIzYmkF92CTmh+HsXUPh61uMSV6pRevbVmayKE0BAYfJFF2JyonAJh65zd
yYWktZbI0HjcOmQ4ExiP6BwAlOskTuJNr2lLtQpR8UgjdtczKVNMCyAlA8GUzlv0
BO7AjS97Cvfl30ZcKv+I78tSIPG12VAy+3l/KgEevRX5K07OlAhz3gSLvkNwyydE
Uw/E03EflpLdbRfKLjtB7fw5tfAA+2k5MOYIqFH5bqMOYmNbhLWckniYLL43c6Lo
oliUeCKgvSpmmd2AApVpGFYqQzgTbF5Tcm9AroM5auzR2ghBT/dyE6/A5uE9eatB
kU4BrS+jlvDqBXHPtvc1JSUKS2x2Xy2vBYxAmUcLLC5Ovc7JT3tnOqKSDWkFS6vw
VUfrRjURvsAEFNSvuRS0eyZkob7wHlw+61KYV3Toyg9JU3WEIkswk0h+6P7sUs6r
MHy+KjsE3O0YNoIy5htzs48SmCRUE5zPSSLAJJSyjk2g6PxVzDHg/unA8jztg5gx
v9FmBibXNOJs7kWpCkJMxpOME/TSnxpeBijPg74AW+ppr/A+aV0R0H3yFa07/5Pi
TvzKvd8PAxZLxrTKghf0PPKrxqYEUCNfQloj79E5ISkmh0XmlFqB7TMcySuKVNKF
fYN4FAO68OU7yWUpxiMO7DuNmhltHeO/gO8AS1gDaTjy0ndY/FsXfNwNmtITRxOW
sSycHy+2cm7RpEtmq7arUppaoRp9Hu0ullxRNYjR5gmrFUaWgS635Qegl2vy9KK3
qyjQEYAA/LMm6eUgmHuoS5L8zFF38F/O1EKuvuTnT7s2IIGoFUI1P0gHXAu3VeV+
GmuN1sx5B4QpR9Bkr9JlQG4kgCTPlF4efLFV+y5jyesh4kjPmGGYlG/s4i7WvOBs
gYhMtVbRr3HY2YDvM2UUbHs5bwDyQ1vz9LtI/2GfKN48W9mTYWlmCVbrDODy9VA1
D+pb5OmhVHcr6jF0PkG7jULIA02335JMe67Mr1nt/nXBJn4RLWgqA6D78K8D5aun
4zRJQ2pvThdtvIwkwaXmlHp3h3NMjblD+EmqKMKme6oLHHjS2OrH883vHu0YQH6r
ldMWoIyCZ04ITsNrJu56TcMhc3kqNguEpQi/o3AjkOJEPNtdS6im7mAjtZB/A5wn
zTlGkqIkeL8OmFVzrYqeEezWxzDPRV6t9y1YDBYhisMZMdhsxNwf9+dHUppQHW9V
Njd3A6LoqrvZTy4CcP4J2OlMcac60ILASkvxxUxJojq5pTytAa2wbQ6wpjUKwen6
i6cglCFHiuoCZ6vnV+taBSWV7tOMtHDCcHtdF3tZJy+u0p6xaRStq8L9ju59C4Jx
ucjUqUKQwZ+ro6rFYaxD5EuxHZylgtn3ndVSAyeyBAcUJypGpb2BhFcRmGXYJSN5
jTaR0JB75jsV0Z6yN8xKBLcNrvQ3+R0e0SeEaWne+1e6EjG1leogtxhzxO+qTE8a
dx8cl8nr0uf7nc1EJsljLXb7uD6UxcNHeo4KqWzk5UcGFe6RrlUl0jAFZ8K5B5NX
IiLvLbpnhUDkYTv8k5zLQWz6mYd8FUoOeQib9ikeQAGoFTt8RHNZjNWBG5FbffZ9
/Vhtw7xPzUbkG2uUwucPNBHKD9zxp1P6PqJzRWXrhgDL6coenZeMdwwFu8pikc67
COpf7Y2RhIbs6WNKJBpchzbeZ7iF/JZWaPmsaVgcerUsnvFp/Za07Zt+RmIDE/9V
MhXDEg4taIKFSTnHKKx0WKV9S0nFJymj1OOEQmXfAMK2+DRAgCSGrqRYrWMciqR8
+VP24wHYVmJKUppHLDw1sqCWD5TTqRfLnS/+emWrQsJiWU3gFlo+tP8PUq7vN2Y/
J+YqEF9PBDUZuIOZ4p0WOcW6qNBg/frz+Ysxo+ontCDFscmTpmaCQoI///u9ASXq
0Aveye2zq5JoWsj1hEZIBgX/sO0Lv2se+wlDHwiAz0WZbgyDdVZC1bQwKBO0Do8v
NAT3u1SGXVVdZUpR1VcUdwuRId/cajnrViifkKNdd59fq6UKfzttuM/au5ewhY9K
TkMcneK2LjatmNcyqDSLbV+DiWlQ4XAPDLVpn5MsFv8livfQ86KhmHrlFWqWD9fh
3eYRJFCDisEEOF/m+9ol7Ou87oQElpvQxjc9wnrZzC+AXnsU8J18atjE8G9Kv3um
QT/qQqfpaXpzU2XAFcYDCJKe72cWLvrzyNvHJA6VuzVbQyy3YhL8Mwg5qbx6pHYf
nCTVHBgRk+U6ZRKRLhKqp2JWyJmAPzY9Id0KqNAElSN29yxdaU6zs0pRzwuBbjZC
+AFnRJ9FpDLrO0Iavyns+iYmtOLnBn/SCKsZYTu0T8xxMzDK1U2fqBNJsaodrhj5
pbKjVwSBk1KwOtlfNk4c2tyoymH0vgfOVfR5syGtuefnyGkVcxt1en6nDlng4dSR
hV9uYn10EyTdg0Cdg8dfB4ofY4zGmPw6MEjXD9iPLHlGsRAzZILiCMjtMsOw0MfC
yynqiz9z4wxHge+7ih7ozF4knQAGibbHLpdfoO3mHI/2E6nnkyFo1QMbEF7P+V3v
pfoaJ0IHQh2F9lTM0qg2XrUuWOPGquHn4LMQM90qN6yDghyPmUETv9OL9unWeyJu
Pi5hzoLB3e3qabX9KPVh6KhAB3lws7ZHr7QknlsUN9QMD+Uy9h8VwkvLnlqxiaHN
OtzCY6n/K9TvpL08fLCXP9LMT1fFqEmeC7wFUjTTb9h8xRT+0jjCeIpvKiGcjrOT
+787sKIml++8bclmfn/YS5bIiT/OYNZtJ1eNAZJU3OUkQiPNeAYLIqiCfdkhUrXh
uIiTt4GJgBfHyylx0mW2zsq5IsgdTOOoezPcIY+1JfdAe/bF7IkrTfOGw0Nw9F1p
8WCCgoqpFzHZgEyr4N2S/3D2omLunqIK6F5cMktWS/1wMTNowl6MsV0EwFohy4w7
3FsluspmjLqk7xP60iegZZxHSGK0RhEvnKc6FzfSlCJrWG3HD6eo//7v1WvsGGMJ
Wcg2y74AApCYubj0Gq/5gX7KL5E3wi6Km/aQWsMcjedSXKeRKw0GkwJiVBxB/QsY
Cq47NwrXn4YLuGgZn76YKsR4TVso2ncJ5PTfSK6FdjMlqjbo2bjZj7GFGrsNu4fW
Q1xdmIJ1xUnFa/mEr43jwBPFQvMCLzc92pl15y69t+LGIXXPftlkgClmJ2LQfNm/
/SqCO7ggdbE7yqEZQv9Jjjf4AUfibT1OduAs7FLfbpxaB33mlkdKCp84jYI9BjwK
V9WdqRO9sWK5JuKmWcxrYHhTp+qkdXP0G3iAo9GCJVAErRsLP3AY/tARDHIGi+Jd
mrhOjfx1/3kKNsxA1+9xiTRIMHO67K2dzB6Y2Mr6oaxmawU3ex8R6bSnhDKp4MZU
I1vWJOM3CLGSxwcGTGnty28DhanTRkylzal1oX5UJZutXVVv+8ELplrwdFU/VzWu
O4Wb8PoGhD9IhB/Zjxgad6iaPL9LrZceIVdaI3UWZlvYR72qqwfLvE6fJl85QsGM
tLN5925vtf8krqFneINk2b3v1nu+r3uFBN0u83qt9uBe8/QmjmtbtqT6c1mAUnnW
dqUukwQU2rGonCoC2G8tGTXg/a9grWFr+SC66zlIILe30vmXU4WkeWsM3qfntQkw
1WNwjlov6lU247M3cCImrBWy2lOSMVw3W0iStE7BZ9MgyjLdp72/8Uq9yDomPGOC
fCqiA8CEd6nnBKNMlMl/8GR4YdocFqfjJFiO9Gxdzrs3lx7zPCxi6ONd0MxNqLpp
HG9dtk7W5ujWBEr1vbWUgB+Cpb+9N8HXhmxBvl1S6mKNJRKqUTeO/pk9bC3TuriW
UCtqwGwPCI6C8B9xpdnVf6W3q/rAWNQHVR2gA6UObjlu+4viAOFw5NDxBiXjVMEJ
y8VpTkLUYMHyH6TigERL6zQ0NlT/uumLd9EYfAY0qwI680nr2PfI9CdZQV0xwLir
vapR8l2swzlejnQBAZB/TjeweyMVG+tAXcMBc6WBz2/MwLdiAu6QMgQSSIvcimIM
3PdBKV3MAnhpYm6Zwvjvw7O2gZQQr2wVlkaaJRZqCahAaVqr8cX4CZ7ypr7aRJlP
p7AFC/P5IvDbBsQUPAp8fMldgCT6KwS7IcNVs4UwBUpcYMP6umDIDnA4JyCAsbRf
A9oePvNlHd9OnvhehFJ1kuJOLaBbszpcHW5kKIkeKljLhqu8gx7YGxOc24J6KrcS
w6RRtQ8tlLcnGAvFMZXEfFHACZE5RtnPHTvIx9cKVG6rJ4x0QrrjhWbcH0TwkvVF
3kd9qnHa+gDC/YZt2dCsfsDaQ7Fyy8yIAlPHDv0TAcVw8nPkpZLfYgwjorvRm2EV
B+58YyslN4C7qsAdogK9i8YdVGFN06gCGwL3u23EAmGFqodF9Ur+kLZA/1ERdT3H
ujo2EjSUJzriu4lV6+RYNMTE3OBwveg44iNS8+oL1SeoltAg2ty5Woi1iDVH9R3c
F0jCxhAyoq2EysgCn7z4YTwFg+xUtkEPyxK6tPv2dUIzfFNBvhDIdbJP8IFCFiKi
ftCSWouVKiJ/CzD6iy1+7dpH6HF35jKrtEkPa9BBnKO2VH/MBQkjy4KUJSfjDfG4
W9yn1aYehIo83IOae6V+Gp3yz3yV3ogXfBeOivMG5PEy25OaXlwgUyOFioEdf6SX
8g90JV1o9UJje2dYVGYnBMZyDbvbVB2a71ULqIBly+PTG86A94pnBsew0DorUZZf
UIhz3axjxH06I1maRVINnlImAbU4rj+g1DzuM2F3GCyQOXMPpbsGDxSJETtY0oIn
fwjY9ruxLJRb0nSBxEGmBvRKHnSAgltsjAyaGZ9SQPdJmhv3qewKuG57UuYj333V
R37VVs6kDUiS+JefG/oq89uMXAjdtr85TBkwoP8mcihhstqO8YZ49yOn9lsp22Zd
seQiqL+4mCCwqQuw4qMT0+5wi9BxLFN9IAFTHZyZctbsB+6vUNRyET4WUTzYKwlN
x7jS8qWD6LJgbGnM3SFRLd4zQOXySBMzYlBHavxizhz9ohgtmxTA2ECzlLOuZO0D
YZtbnrDpCgLHVJY5JgpuSHLbs3PkJNYjMlPgRLaWqJRe6vcMYMCJJmQ2kKM1ZZLW
d2j4DUFYcRNHXC846qpNcg0JGX0Q0i3s3Qd5O+kh1gHsCVJh7lHAHgar8aRjsSKE
FXnVLDNAapmEhQjQXvXSA0tSSqLkdv279lja38B6ERlyWHHMqxYhKDMXAXu93JHp
HDSlZLrv3DX6eIVndsoLTerof2NSRoWrY3b6HkNRs4qHSvSkWIdaXNCsb7UBYDjR
XugGatTfPU9Vp8/E77cX/2SDgOjccSVMdaVfaHBNOQ4G8bKMhyKVIE2aEjTLmU15
KZC7ne4uiRSf+OdzgMkOTgmbr3djVg1zuj9RSHrZCYg7HhK5uh3tXkxoG1wgKyOP
ALrQcatAe8mIq9uVrJ/KPhpDjDT6Gw1zPrmSE64aHX0XdABNnRmIg9O0TiCpRu7y
WqO+r+i0C/Q+egUe5l/mmcfH/+bGc6O9k+HT1EMe3uK0SuwkuXWRGNrdQ+PBQFi0
uN24Pv/uS9n3IMW5DF1myRIMos2Ds776CWr6SLss+lLXEahjD5Mi05mWHm0sdSB/
BeP2Hdo2VwD0nUcuSaDTWynPcrP9tX4z2R4TxtpYnn/mdsDnOGkbyCW3XAoqu4im
iWarcue3L+pN9j6FfxWArxL6cJgrFE8Ic0xEDgXHU+emPFjqtvMne62mNrFXW1xx
+tRs22A+kUFkz+xFVuxe4ZvO83j3Yz6pRicnyDCXADM283PNUlvY/nom3EAXyfiA
Q15YPXlNEEgeMRGfx5TbQQyHgUx0jaH9SJB2252KC54jDmJeMtQjWRO+CAg+Q8Wj
5O52d3qA9ikOUoyDkT5wExZyOoUYYQG9KXZ3S0rNoHgv/HOksDRUrhBC0GsEsMhB
p+eVTNioJVGvqfURD8qx9mV4wd1QGP797ARHLVCofxjpoMqwcgp/GpupNWdlpQeL
v0Z78heYayHYtgjJqeGaDCyUPJV8Wg8CTLgLvllqi0MtPoRndPLRl0dItMXv96YN
63CIqWIjG8Hzm4cnB9bjaZj7y960TppPeo8BMx6FxqbJap+LV11namTEHt12hyP6
nsfhfLJV9G6yMK1m363P7GDgYbf5GbFHjc+RhDroAc8WQRVDmZSalhb6u47p7kfE
RK/6Zsi3MJYrsKMiPqRJnDRDsalS22mx07iUo2QTEx1Qi3AxTq2UU2vYrIpi7anP
IuTgcdjazQkLTlVdScLiulpNO521y7twbibyph0isRDVuQJxIdls7VkALqMWTBjI
Lf9IpaDYyO0SwvDvDsI9WedxnAO+iu0jJ12xo2A31Jt7JODHSnMOj99IXOhaakYn
jIGzb9ZZm/+b1v8gdPhYMGwGGlz0FbBBxPDkLlnYwTIZsE+Nza8QsZ0Md+LZuYTF
H8+KCrikStc37sgqcRNs7+2Qc8aZUAvOdSALP8EHWnTSzynFRQP9ktIJbMp3KcdP
BGFEjBHk0IKqmxbcXz+/2jrW4nY8aNbdHROljG+6ntTUyhtgCp+esBhMFIvSP3n2
g62YFrXTYVHbOUTsNIDsjinolUW5HOGQvm8lRdLmRq0FpzAcxa6znrKQAj4vXAl1
pf9NqLWRg05lDOHLHo5gLmVcMlwdpOeBchlsl6Ya5BPxtu7EAS12oGiA6CbDmoeX
rsOYuOi3rHJR60RWLiw5vD3pyJjFb98qABgZsvbjXhn0Flj09xF+IsQlney/Fdi9
3/26b1+mGEq+aeibndb3bUc4buf2bsMsyJsRwP8w++mifJmZt7FehVFUe+xrPKOe
ewJzjKC5ikD0gUWc+wDfYmw3bQaBKGeXElFv3OTDhdcdfqyglTqa/aLGyFzUZp6c
mxB7Ay0nhtuwp5SB8cujlZDXFvL4KkNsQw+XqhUwaFNKhVFytwYuoaesf1EOim/i
rhdDyZeP7W6sClJa/1dXjmWm0FF7YPP6PBsLdU45g2kbNg3SxhhUBTPk9MVF0TWP
QXVCGxMPYeilRpQzkCPgLB/zrrQr93kTNEG9AKqaoR8WpvOLZYacNScVs9PaggLE
ZaHB5/gJtIW/bS2ZVz1RdFcyd/YFAkE4DaIMIQkK72tlJeW0igtRKB6Yr3pR302z
VWjp5NZ+MC8wwrx/ccTMAln7XPkUvh/8b41Pz9xQS6BzGS+A9TV+/VfQ+rB8eIsV
mabLuwCpgnc5nKVJo8x0VUIfRCUB2L0umX/Wmb4uVyG/71ZFUL/gZpLyAEwejErj
GnxGoOZoBKUXfkCXQZ2UZyVDDe1xDMFevCDsY3KfyNPjRN98icR9zAyTDMGpNWJF
19E/n0CWpZ2cgSF+xtWjttW1WOR+V3iUCxeqZOOZKv3fXlZJ8GYOARX7V+74dAoY
pD1aBFSFYbMqSL/rzVOI49qghqUgbmI9pQrZhOuLEiPPUFSFGWVZhagXWLEXH0nx
ybau+ijJfhkcALtB9LB8UpbItfJObxpc610Qo7QFkgf4/QYgReYT/6Dzo5f09SUD
v7HKvcc9Won9CYfRahiaoxsxEztA+xo2qKeklmU+1cm+WOxiz/mY/H4zzsV44EEU
QfcPE6aRXUyxUSn0RqR62g9g1YrXKCFzVAWgTIstNX4FBoJ0DYfnf2Q/gYikpkwr
V4SJDpgc2H2r5Zp0hGGOhgrkbOmV9cn09sh+Z5jTantbcexeIR33Wsl2f4He+CfR
E+Y8tLb/hGDRn3VxlyCOD5TxqICMA0i9P2kICDKGTaKw7ymF/0ZzUf3vvkWUH7Mq
IjzbGrwD9rkmVa0059zGrD9xPYt/kcYSKFSGlNs7ygNemXFtMaGEy2K4VH3mQpag
4poETRuRj9sQUHwQ8UMpEt9pHTU+98iIsW7WQ+wvVw4e+GJDeiSjthHlQigSGAXy
7nALbMYrnpqPfO/ZE8v6xmqUYVdxH531HLWH+ECrg3c4waz8p92twzIr7i92Ted+
jNhzjalicY+o8QHPrKPk66+RS2xGI40DRGeEMUM1eAPvN7gcUBOOJAiUXjnODKMk
2cABtn2HoZc63ZRm8d/mou4OtEdbleJcjV6LXSZMsCuWvtuE+hGkM8twxudzec+Y
jQXqY4J+/eN8wYxBT8uBkISwbNvLONsphv6uZooNFscydTjT43OU5175zsXe7gPT
/W4GgfZ6zNIDdjemPHSNLASHVQ1vT+9CmiwaJzi7lSC2P/pn8D46AIittDKunX29
wJuUctO3EcDJH0ooSmZy59mQd03SvFyHJOa9abrkYToCuu+sffw9sonMvOizvLDU
MM8jGcTRZ0Lvo2FpoIvFGb20DBd01hBxG4xARIqm9RsSSC1uA9YtYhFjYqrGYV+k
oEIilwsJjazWPo/7SqZvnXaGk0U17W/pBx+MtagOSPZ4DeRrfjaZcq8HfwI8tqbx
oy0cUoeP8Zlqbn5iIMIVc0d4WvjIiTqeC4sllwR8FT61ztTrlf/7RR/Gd1T1hkZc
dZpwMyARGOkQW3aV4kXidHFpFu11ynJbZgqDRkoNciLF/uD6co19UV5Y8+MG2d2X
s/RzebpizX9jmgG/NEKeRQbXMzPgmGnw/8kkX6D8DbCUtZof9ErlQwHUeXLTTzds
XwC8B4srxegnS2jzxaGx5C3PFOmHzOa2jbci9zB/yOcQ0Usj9IHha9yO5UX+9IYc
pgCDG/zD1vdRCam4uBaE1k5I52rckLnCNP67T9s9VUPhH6TxbyPAinp1U0fkdQrt
T2NKgh+eJScSZznjVEFJnI8ALfbwmDjdwF2zTHlB5jIDXm6eYE8j5mOtoHwhCBXe
8bI6IF+12vTzVfK1wXu23MNdzHLr8LVfSGb7IQA+SiMEzdZB7RAUiu8FldHRyJpC
w6JKgw25HhM54OiWYn/PMfpb2zXzHB+OPu8mXPqU0WhB0IbflpJzuaP4VCTTUEWk
3swfsDZcrRZn7JR/PKJaCOI5y8+j9WrAreI3YXK9FyMpPxjhna85paFa2kR/Axrr
mW3+lhHQQmjQsC/+Mu7dR5MLOpOZehUunEK4pbq+wENKyYBauu8ZE4aEcsGTWuL4
Ey5nC1ivZjOmcntfi9/wMBc95HNDavjJYz5BT+EcKpS/suZ231IkjxKm7WtX1lNY
9KggizkZz3NKHAhGGuN/zTw2DyLUZ6T/t6JT6o006cu+Cdi5szZQjAQ7/pbNQKe/
cWiVLkxejky4GuerXUllVmtx1GB7NSU6qvCs0NK+fLAAHaiCwmQ4KNzcAHRDaeNE
ZEjeHq0MPv3zrjxj7RDM5QA0McYP1ncdIjPFJ8l/OeaOuBhp0Tybf8Rh+NnLtuiN
KHgo8AI1fRUYNyDEfFth40A+jf0wN5DIUerkiUN29Z28wkcpkT4CZmA6sI/4Ja/B
bSoaM5JaTeuVOXRUEDwtBBkvS/uReYcwGkG0sHoNr6ox7gME44h8IugNBIxpWmcP
Zo5mrtPYZ0Qxp4Y8OBI1uGq9P/fLkjKoVSByP+YwTG813CqHgDuJ/duMcDMYNa24
BeRc+G262to0BTk6JUd83xN10LNx1n5+REEJipjgvn3/IBU7yU/elClaF1nY9Sfx
FBw5RRGQm1+WP6NepM9LTmR9UoJ7NCpFhRnbcwEBlsTCZeFzx1gOO+sOW2x2fRzv
A5IijhOUowQA5vOdWCs6vEREz8fdMxkgjhN3yqRbMmvEcBz65KAbUNdjVn6NOxTg
y+GOzO/1PltdNHwRWFlfpXxF17EbFhC0Y2aNTVi2Gp7NrOzaqZZx57tA7yb6ewVI
0GlF7PbWy+9UYomUvTR9ygVMF1pVh/lP3nhMGNbSnq7UFetsZ75/86byU0rco4ia
YpN79Z8mZI83JycbSS/uVg==
`pragma protect end_protected
