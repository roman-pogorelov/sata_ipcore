// megafunction wizard: %Stratix V Transceiver PLL v17.1%
// GENERATION: XML
// sv_sata_atxpll_core.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module sv_sata_atxpll_core (
		input  wire        pll_powerdown,      //      pll_powerdown.pll_powerdown
		input  wire [0:0]  pll_refclk,         //         pll_refclk.pll_refclk
		input  wire        pll_fbclk,          //          pll_fbclk.pll_fbclk
		output wire        pll_clkout,         //         pll_clkout.pll_clkout
		output wire        pll_locked,         //         pll_locked.pll_locked
		input  wire [69:0] reconfig_to_xcvr,   //   reconfig_to_xcvr.reconfig_to_xcvr
		output wire [45:0] reconfig_from_xcvr  // reconfig_from_xcvr.reconfig_from_xcvr
	);

	wire    sv_sata_atxpll_core_inst_outclk; // port fragment
	wire    sv_sata_atxpll_core_inst_locked; // port fragment

	sv_xcvr_plls #(
		.plls                                 (1),
		.pll_type                             ("ATX"),
		.pll_reconfig                         (0),
		.refclks                              (1),
		.reference_clock_frequency            ("150.0 MHz"),
		.reference_clock_select               ("0"),
		.output_clock_datarate                ("6000 Mbps"),
		.output_clock_frequency               ("0 ps"),
		.feedback_clk                         ("internal"),
		.sim_additional_refclk_cycles_to_lock (0),
		.duty_cycle                           (50),
		.phase_shift                          ("0 ps"),
		.enable_hclk                          ("0"),
		.enable_avmm                          (1),
		.use_generic_pll                      (0),
		.att_mode                             (0),
		.enable_mux                           (1)
	) sv_sata_atxpll_core_inst (
		.rst                (pll_powerdown),                   //      pll_powerdown.pll_powerdown
		.refclk             (pll_refclk[0]),                   //         pll_refclk.pll_refclk
		.fbclk              (pll_fbclk),                       //          pll_fbclk.pll_fbclk
		.outclk             (sv_sata_atxpll_core_inst_outclk), //         pll_clkout.pll_clkout
		.locked             (sv_sata_atxpll_core_inst_locked), //         pll_locked.pll_locked
		.reconfig_to_xcvr   (reconfig_to_xcvr),                //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr (reconfig_from_xcvr),              // reconfig_from_xcvr.reconfig_from_xcvr
		.pll_fb_sw          (1'b0),                            //        (terminated)
		.fboutclk           (),                                //        (terminated)
		.hclk               ()                                 //        (terminated)
	);

	assign pll_clkout = { sv_sata_atxpll_core_inst_outclk };

	assign pll_locked = { sv_sata_atxpll_core_inst_locked };

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_pll_sv" version="17.1" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="pll_reconfig" value="0" />
// Retrieval info: 	<generic name="refclks" value="1" />
// Retrieval info: 	<generic name="feedback_clk" value="internal" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="ATX" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="6000 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="150.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
// Retrieval info: </instance>
// IPFS_FILES : sv_sata_atxpll_core.vo
// RELATED_FILES: sv_sata_atxpll_core.v, altera_xcvr_functions.sv, sv_xcvr_h.sv, sv_xcvr_plls.sv, sv_reconfig_bundle_to_xcvr.sv, sv_xcvr_avmm_csr.sv, alt_xcvr_resync.sv
