// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:01:49 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ALC5o42OETN2ZVkojUcsL1ahPykuuWse+BurZ8IJbsGaOJlTdTkMZ/bQRP7ARWzJ
rA+/RyqvdxRfkJXlflp6O/xRkXggEQO0YL3O/t+/VuU3FjvHlQyTW/QVWvAvNgOu
Xyqn2FruKVjcy9FZ+49Bg3me9OZByGKkoyl4tPTlxEc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
ot3vAJiELH5uB0+0/+06v1Q51z++kIvSJTb55ro/qVfmzPOp6Z2fb/wW7xPJqz8Z
nAGO5gd95JbDUG/bbw4XiLjY1eKDJi29E/R5dcSvpUIib21WZBPkkkso3oxBHyCC
FqJXkK7UgSOJ6Du9RnkSMCZvu2goA14feLYy+Ck8j8SOP6rr/DXYORcDtK6h/DtJ
5FH0TBCV4qiYIgSOK79cE6isjgVzUskv1sDqNmU//rZxc+h6MdDf0ssH0th4NI1c
+a+kE+dwV58kXkKAw4XHUcaLhcskQd8KWSxuAtcH3qt/Pzl8LzMdKOOZeCsOdjzx
kC0b/JTZlbNOFExhM8Wm2v7XN+VLNs0VNqj68EbSoe9bCHf/ACsNyJdThjqX7FWG
DT2WFU6PgQP2Cp+0hHIvoj6Hs6ofDNMVNECRZT1rPOFBjFUNhpl5dpAAKWFqnL3/
ZBSFfUtDivuX8R5Uz+tlIaCjf6fzq9AV0yKj3m9of8kHW88a3eo9OMoDhgSpz0a4
3S+Rf+TWj+E5VpvCMevuAInfy7/hf/j10XzvYPss7UwqwAi+0bN73M0s2T/QMDNe
5X7vxpLKqO5KWGyre4n5dfGxtOYqJ+BRIm6Y1wGNKAQpdKpNfQG+4avm9c16GcWe
w1SuqZRr17oJnlv7V5MNmmPlN2pRpQqf+WOw+d89gOuHPCQNSycML7mUHM5FUPEQ
4M9qh+uYRjnAMz91Mb+tGF+v7XJ9GeqGBprLhk8dFiK+OX0YEKrC28cspbnsdco3
1svfkDkdUJkTrHFnQAF7Ibea4JMJnIztDC5W3SpvR7LWXbMmR32l+bP2X5KYWJn9
v8Xukoe9W3jMRWlmpwY+jCoejyrTrY+lZiERZVx6e2lgg/kzUuEzz86VRThc1jmn
x60usSXO7kHLi7cYsNkS+gOYmFZG8ndyB0EtNJDwqZt3ngc5OK2i9ttZFCT0PKgB
/Hbk5N04+U1ATBxYNaN5+/1myP9WWkRcPPQM1+9C0J3bHW71Lf1VeaBtTMl9YDcI
C6fF/Jmhz29Nfqi1o/wf8oiPczN3v7nw2MmIDXdCM2k2EZUObaWTry8609vAmluo
E/Lh5e7sC2q98NBL8HzBUb7iEG+eMBm8wZchinYRqyJGdJyqoF96+2/gfyuJARRL
yva22/UKOKG7T3eU0iCVwV9tfPBWazFBhiLJ24LvGcpyvuZ1wgIZn1+zBx51sy8W
YhVtCruniRr002b8WRFH8XzDe2NlOy70xogI2P9A4utukdzzHongQ1yGxm/DiBXD
05oSVC1nD0UglMnJBEXvFg5s3U1Klcew8fYwUTWxArk43DrsLUY5Op2zKDJEnyOQ
ApPBPHPiuK99mrfGzAX7xYO+yh7lbvLQuwRkWDHNEqhNEnR2OItKyfwCMtUusfGw
zmKgoHL/T0zgkPzm5X4xrCjq7FX/Z++QbiGXtqrbQhA+cu22hDHP6JRzxyNepqgf
/sf4s598Cjnm5VZK/ziDhYg3BVy8rqn2nzzu8x5YF95SHHMaKaQlHmj+YDHSrp06
efNWAf7Js553x4h+nDRqsmJu5QuzHv2S1ENQyo7xH+/GGn6hWYa63SWsN3BNhwY1
wvcRjLauo7e3r5U8Eibch8kediBfvIqg8CJrmvt1PfmN+TBXKcg96snczkFUXaJy
imblawP7KCKIBBusjtltwyidQIwj0naIk8796L6Efbw6JT5mMStOoivaxsC+qafc
6MQnPGUXRxBFRoUSMLoDF3HHIk38/LUoFI70L7u6xGhjn0L10+v0A2xpj0efgxcY
rBW3LPvprP8STxTfLB8CirzEK+rY9nakPk8k46x6jAA5tN9yUcXqU0R/RGlrRV4G
q2hhM90JED7i6Lod7n3tpkwtDMx5uN012kcjLQ1CfS2NVeB+YjmHsWG8yAhlAwty
YJhSIAtUnfrDSohighVt0XB/4StseeOz7+Tr2HurdY/WWTMgrpJGRIsOz7h9kv3G
wzDydW33fHEtHq0D5cRpq/vGVq/seJ5HaVQAmPbjNTXSoYJIdKcXNeBgNQuQZSJY
eipJa8MA9G23KhRthUSH3Bx/XcCTUsew3msZ3NfijdWdNMBtUkQUDkcigxTa3TGx
B/DwFNmrm82pKxxqOVKbnNkF7LyPdWpVBhQVH7xNTgzLItoVJIEY3E/SUXw/Kdq9
gR5McDNCKgefrUkmq5xNOZ9yllzzv6KQsbjFKGTfLLErI6SSk5FDhs84nosCAVWc
pflSLEitW5enCyBP5NCO5phYCtBdZ9si1eBBFqWaR2MuhHoN4mDKBWfLyTymWpse
XxnzxevHOOHEDv2Bh+ohhF6QqsOMWFLnde9TxrPojUnu9qcqerUneNn93Cuobm0h
zlOLB13y/LPtz88j18leOaFuQYUsWVn31I4ehHMfd6AepljlSGJq+s8pFLLw44Y+
lRc4/0vXDpCKuJeiIOT3oNR9vJiNGuyWUqxsFgqz84twkw5+KFetmwOwmbLv1w1E
Ip0efLvZnNk8acCno2f9F9j61FDvTBYt4HmlajzNqz9f0iAw3Tmqz7Rf12J0VIPS
Cr03T7D/cXwj/yHvJMHSjqwBweiAAQC1UJSlg6GRWFnPBuujwYry7cEN5gUqcuxB
4u7rMUqw934BrcyhGzi0sQetBFE6VJGuBD5b0ORJLNd+5pABKIrhf0SKWYlzH1pT
sFzJNTv6PZ1izBmloIcyNsQjcyXGaXcGSBI42yVgjEwly7W0w3ANfLzY2TCYjI48
llaV0ich9XQL82c1H4xdjiGIS0GseMvhmTAb/8zdMUCNj3rS23CiOu6auHq79Ikk
hK/smnqHC6eyhSW36CRjTddL1nI4CPleTZbGVM4NQGd5Ix+MXSFh75ru9Q8F4bGu
dpkWrfzI6baf1HXsBVOpE/5CLLjPv5HXwAm1fQa1+M09JOrfxdot4mP0DWpcSDcq
hlG5A5qf8+xkGfdmvokIduMaTbr67bv2kffspIynzX2zjbTImDNXWaquxL0JcNUP
1RPY3GMVj6xKyF1pqX1P5tc37Uapcb4fExFRf/k608Z69fOS6t0NYxfDWAXqU7Tp
mjz/d2yWdRpfrrO4EpXRyT1o78CXL+wMQK8/+yW2DtsFCAVCLiaa12hpAE8054mu
EGDzAp1q4RIM1vxdGlCj2W+9gvXpRbw0T7YNMdoLGMtYKI0j+pbPw0K1vg1A7/kU
+PmWgXNKLsHspJQ+Q8THpVV6BHbz28hJk+WQIlkUGUxhvFmQOARBOseH9c8iYCpP
qAFCivSMOqbWv8GKto3dk7VTDjEHE/ux40zpAeBf8KF/y33I7xEgLsyUbkuczigj
2aRvQQi6gBv5pykWrZbe19SIsFQAXY+xUeAX1tezPFZbMY934dPKMuPVj9bCgMzD
tSyiXTREshBRr041MbwY/8QoW4HTsQVyX2dYyQdqb7SdCnX7FsHzXkKFQcEwiy0f
c5zRpo6epzr/I2k/ccRaWDs4SgF3lOeXo85sySz4jb4k7sK4IfodQd/tZFt3gtkT
kR8rTk07uf1mQYDRl4f0ddtXQlY/esjgzoZICkEJB7sxthNtL+Ph+EyLzBnBuzdJ
T44wCfDxVbfn1VcQmEMUunwLSZuNIeFuf2ilfQTCCEMzhUi4oVSRWN7ctZ8M27ML
cBE0QJ3OI/JkTzDlt1sX+KAeuRq82YNSrJc8bxzxkE6gYvLCPyoDU3b8OHOPT9Vv
gFWUVdzDdRl5tqwGHIXTBFjfGkyNX/V898VxSx0zVHqrQnWm/gcB1Nxhv7vOKo50
1yBVoFr2baN1jxjGElginE8kY+HeUMtxISuPlN2Ry4OAzOn+k0jN13MU3W8wL5MZ
oN26NwP8YKtVEKiA/2wM/rGI7g5fFFMUV8l210MZiWOg18Q1mGSHrp6cc7R5Vwoq
RnvaIrPKlOLQcEjQcEeG4Wjh3QCIAaau+tRZwYKYaRBtIOSz/tNBZ9q9epzVUxLi
ITDLxo2Yf5OMoAbRe2pgF7mPOo/btLbNebPWizlxg0ZFABIxdylthW40F7kmsdkc
fyQZxQtCqTYV7pS5QFn7+hFyIQ09pCwCTWRmKKHHyvKsYgJLj5HI3s3flUebwga/
pJsSQe4nVo+DNKNCULhNoVoO6lNSpDa7YA714OH131ntjovdHH0WQPuudpSD+988
PxU2TsEtmYjTzYQkGOhBQhHwGsWPLe2ByLJ56SHKQ2BYBCqk6ERfaQR+twNBNFD5
6WM2vveyLVdx6PDM0MFB/79zBT3H+S/hp3R77DQBxBxiMvLeFo1GHQizMqwvGn6e
nYCLtuB9QMskTtvWvsHtkLjGKNViXQjgGShZeYk91d6DJr8KSxv+qQoSpKCSWUTv
wouy5svX2j9ECtaFbFUBp/S+WupyYYZ2rz/YIvEhnXbLH9Lz175IzY5UBfyTKPrg
UNPRm4KmcscSw8ftFhrsryUXsLPRxemHh3lKczvO1se1Bq5GsnfzAVNZv5oKLoYD
qjCp/1p8XTe/kge1EM5b1R5/b5/qEqeAkn8zhgBkPThTqxdH9pA41zjqjVS6icID
Pv4Bm9IUDrbczgIO1ZS3Wi9uvkT8N1OMz1yMz3ge5RyFWVAtkhi2IIMwIlnWItqV
T0sOoohofou/szNDfPYGIbbpZQKkUK06u6ZX1lPuusiV4jxVkPWn9Symp0IsmoCT
4lUGvUiUWY9hOqRKe9Xcsjyj6eoatUKQx3/iId8ev9JDI5cX4F9z/8yXFpRP5Sk7
RHUDGaTiv3Ejs/3aFkL9XIIqGWCvuEQnVfaB42MVb9oyVALufAo56nVCOHCQH1W2
kHTDvpkYZwWUWygTSnj7xCWzfCxZoukJdkP8/GnDd7Pc53+wF3xfSXEJ/xvesmTh
qsdi1+q/x3HEO2hb0EOAvYtImy7daJAy/O6iXkf0RFn1df+yAKZmQJQu0+RyX+DB
H+inC/ZO9487U8Y/j3V3U1fsv7tOEycktXeTL63WP4dLqBjI3jAUqum4NApRNCOR
5QzTy9PSSUMey5umzVUD0W0fPx4AhMeBjA6OSTpGs7plYO5blM1KoLC/9BusqF6U
CHVeflzgveHkn+j6OIjf36V36+67X07otyiWPHLfaS1dMQ27/Qt9dF+F9KkOOkL0
86y+K+QRjoLsFYdyGHcxqsNIKzDc+SM6FJAsIIlkSNbo+LDpUqkKYHqNITIvqNOH
v4ccun6DpBBCOc8fq9xEX7q9HNwTk8iu7GRYr10FobRN2/E4df9CGdz0/WDsJ7IO
MIms9LgyGruwRCYBsCvkTt6Q8QfBzKG7CaCN69ORZaKa6zvwVlnenyouf2coFGmF
zr0QKiloJyyPwFN/mnxAcXf/39R8VMkPF/26t2FAxUzGeuSlUBn/oF/RQoVZZXBZ
8TKW3b4id91EkJaoYuLhFGshQTkqBKdTLNWkoHFRGiy6PlvQIm6z2VQsltZvUcTR
cnDJFTvKdMV2B/Koy6znsqKejGAssYPSQZpwvEVB1bQ5No0Hl+g9I31Jl9iYcJdk
dqFZXk+EyJFuaIZB/hg0rtIXVEzhrDGxwVXDCmAsaAlymDDsm6ApefsmUE0VxDb0
jw+bSAl2X4b40L/bWtsMRChUx3AlxZ+b55yILRllA3fcIs0nhOjVQP1gAzKncgjz
25RcV5AtW5FTs11aK5+qF2FVwvfb4WmcNTk0KNMh6nCxnTF7aqHX3Px5Ng6q1B4L
iJGbRWrYzWm2/W+F5RYl+1QztRPwAYP+dFgCOyGMZZ7ltC0Vdd99hX4UIhjcYcCO
CraP0hov37RemF4AJPhT4Q4XKnT5whTChMIyAsgYSNslZzKPpZXJBNgoVs1ujsfU
G7uVJhVg2GLgmNgtV01CygEOmV0Jb+8Y+cjGJ7NtHf07P13OzwfoMKkRPHOmj1G3
gOxW0D67coFbqG2IvwPRwAn4PGaEzlA844ECVavGSiG4K6lEVYy6CVvnEm+Pd8xT
lCdGmzLInK49UKWqvPZhI/N8WZxSXO+FsPJ0/0R6c9mQMLsPu5+WFB6ePwOSW6Rd
8aLqjjf0aGZ9grxyxqi0NEQ2S5VwXa2WhYXZNMle7lbCDznxvmGepXVSBxCFqu1H
aCDkHhz/LsnQKH5oNDxCtpbTyXVT216uNGrx3CqdsxYZSLe7Pc0TNmAw7Rh4Fbo2
/bCXsY/9yFyIiUVK+wxf2FnE+8ITyEtY+5drpsnS5TFtq5Im+CYUKqI5Wl9lITvs
nB4ulX8QUMjbS0mwd8095pUlaq6uECF2GYLCMWq10fcQPEYaaKOB/MKqD1Fsi5H4
F0NteqS386xnYVe9Z/JAXFSgfLg6OnyhdxyUP3f5HBVj9CUoSdIhDLGXGmvc4MUw
yTE40Wsk/NTpNYU3W6czbU8JAMxRYynRVCOEvKfNMH5sqq08x+o70xoqPBBGNmKm
Drz1d9Iif61HZn+T0sO2VL/x48RDrj3JG7ImYOrvxZs9IVhwVLrkgRCEBwHn4gqU
++PGBlRkFHNApmmTigZ7sPRrJ7dCAltdiooIXAM3llv4c0n1tfxb3duUfIpDxFSB
4mwB+p7SrMG6wXbVx26A92fDBIHk9qF8UVAdVJFF0Q9+O1bgurqLHYPHBGxqVmq0
40HK5ep9uj2H4nlcx1kHajGEqkbzO+KXhFl277YmOei7709/tbzlpeXMGhckeBUZ
p9N46qOiXOiafmRQyTJXabdTElU+h58Nj/j0+hZOble+V/xqh+1Ge2t/fCtSykfH
sMi0KIw0IOUULL350q5QBn3v1rtyP80oT9pH+JFO8QOK7GWRx0nGUy0WH0eEX1AG
/FBwplfrMzAhzVJou9EMHugkkJvHRHnQ4f0h18AbBCuYCwckes802l01Z1Uebw9t
61VbbEehiVF1xjLLMvUL85m9NfGitp/5PTEWr6gnQps3J+gVQb/m586TvybXI4aM
ONNPN0NQBxLIGphPhurm0qlVNLfRkLR7mcrRZEaRuDIOSFZXRFPcQTB2EAphIDKz
y5+8fRiMkRYwvp0ETzqnIH+695znEhneMLVStAaCe8pwBa7YT8WuVbvtckHZhEgc
W/vrx7h17Lid/6Q2uOnejVRtYDrlQiqTwiKwDFtie7yEjTixRCTGLToA22nhhsp7
9f9twt1BuqrDD72YIAs5/WB3U0HmjekmFq6zk4GPV9bRyUtJ9sgwMaG+55jFA0zQ
a7pUPmW015tJY1osYI1sANw+Bcby7uxbc/YZzWDLY5bxJGmITrzB4ILa2XKbeuce
JmBcLb1M97aHDrURud6Wvw+uRomBf49nxK1XMKH1ijhE6J13g44atDL7HuLY+MUv
jiCPOLXGHN2Gk0utHpv+dBKYftmEhxEnS1cYu0uCEhp8wKQRbvakNPL69b1Nxa5F
dui8JzfpO1PlhhWbiTnfhllDwfz8qzVv8MsWc1nhCilHCz0OFsM3VQ06s9XIO76G
82qN2Sx1XjncPoTbDrc9qwU+H/JOLsP+mzKyyjINOdU7c/A9XFDy+ufOQnBRg2EZ
v2N4slXqaqbzXdWHrOJDzT7IyYmpP9CM0LXYi/oFKSnquGPOFq3zHkvEWG6OED2v
Fnu27XpAqQyqtf2XtEj+8QMcPjoORUHtTZOnWJEKSIXFNtqkgZ5mM+ueEzH1KSSM
tl5Bhbrx1COVxHP8FN9KMJL04T0jzhuqZkgGZzjqlaOfjbGtz+D5KKeOvtpUBAya
lNh79XftmD865ILDqIfUM2XZwfD7wUzMKvs7OEv+rrjJmHb/YlgD+Nsf3aTj6rvH
whh9UCsiSPmODyhDSlpDP1CMl5FuCLnkDwKWh9SmibNJBRlrrNMzfTSFnKn4R0At
bYp5h0GcFEVxbyiBKDc9EVsQS5xSOk6CNo+uZkE3bSCXlFa+0iFwEMDZwIAwLnG/
vrO7HIPybG1vxoTOQw1qe/WqGzNuyxb3Digw1H+tY4X+hEW23rS0wb7eL2J5rkCx
RpHEPnfzP975USKvXtl9oyvloloDkd8mPZM9iLiIENyHAi4KTdkgbW/OLK/CSrhB
YhnAbAung+FvAjrEbctkzyyZeMbQke9JOTt0sYNj/KOE3N8dV45ZZ5C4EFoDT83I
ZrIkQQsD/40PZZy5o2HEUYa4eS6sWaFA7yh7+3xK2VaeVHYeNclqIk+bdt18PIPj
ouOO0py6/XI46GrSAfYLAKyeCnYfPoTUc0zsqa325DCf0njFtxVTtU9DTOJukdbn
K++BvutaGTQcIu2a/R8/0+D7OT63J1nfsd2GXxnOirlNc4UTxFxa8hlRcHy8J9Sx
LpHzJlGcDMq1HIxKy7tLQN3jeIfIC8eFdDvez5/NGKRF5y/E+cTThvzdYjG3+tOH
g+shqs+0ZxwUT6AnmnDOnry3z18MhEzs/UwUhYlFN27ZDnLfF+sQPO0jUJ6GRA5m
2HBFeYRQnNKm1dmBKT553oPkaskGs3WGA9N4okVVHtmhN230IsmpdWUH7oGRIWXh
KPyTWGxzjFx72JH/jA172/SK0wc5b0Q+uTDc1RCD47MxCfT3M8tEAOwSS8H12Vq+
UnJlwYNawUK1uctPNZGyPAv+w73C3l5nuDA09ADpSjEYCwIrT6xaMCiBc1NNUYq3
M7FqIHVXg3WdfOVN0iUbI9iY8gvdflCWMRMEp0ccOMysZcHe2twHMKODoXOSAQpN
o1pa1YiD+fsDSmDFEjrRdsh3penpuedn33sLHs8OS4vmuKWMKsGXBvPQ41gouuSb
GmXk4YYyH1gqRX1NptNqA2GOm1FSp2iEtez6cwv70idtHtZila/pY2b+U0aJVKHN
ZXejpOYBqlkkoKL/s8YyEA8TfXd/NEbKFjMpg9D9AOHsWucSElrPmkv86B+Is5xA
8JFR3DL0gMLjuJFTmUgB3kqaglaj95MxWIA4tYSgeVXqR0x1Ny5SaeCw4VWuzBxQ
oOLD2zX97yz++JwWVh45tzFNuBOiqzaiMHbRBnWM/zZApvp1X5jDsf2NssSROi2S
YwP/dqbOKMEOOj2nz/n3NR97zBNgwzHsfaonnFj6agctnqrPbATEho3a1dqfTOh5
rVp95A/8ik6AOcGU530nFC2Wl/dlklLVUxl8OAZjORVHBxPZt7K5J/TDHhpm6s6l
T9nbDHt6geDbcd9nGi1XJKQ9uZGLWeUevrhv5Szc7FnK2KAjKgc1AHhcdtDGH4Uk
660O1J2xDurIQgq7im/rr0IOTRZHxlhtTAlT5YxgPpWzN3/9Zx+glMYUXB3xYjzS
Yf7OjWhaoly2EvgEJI5fRq7yjWvDT1KSEu3MbqNmgJlWaNdJd5roGjAlfhf7tXQa
ZlTCPcHgKmfqCYSIrG5oTBQEBDzAlTJFdCRN84PWMFfMFbwb2i54/kjiQpo+zjBB
Z/KKNImri3d4RTFSbjTAifLY2COkz4nzI4kxiZ2AzH30S10IIj9AmEIeLYw8eAKu
hxi4bWScIWciWKLhvYr9N0nsLcumoIhPO9lImjZtAC+3piBWzzhAI8SFD+u9hoyA
2yhQsFfGk5IzecHVb9HbU8YbaMAg6dUVqG4rBtn+XKwCrHcsjfsrL6k//pZGx9l3
TYnDH0JhQtX060BaeY0qjVMyMlC/GMQMdzeYJOfW4zCWznM6Tr68jlAx2SHMthOs
CP1NIxWNWcYhOJ6M4ckpjRHp5KkwGNbM9YTpECQkKvWJR3u34GE6OLbRj+LxgFJL
5WAwuro7KKIfqR2s0Yiudt7z7+XDw12q56ZMogHjxXt5F69BMr37kOrosZPY8T3e
5iL0XujzqZ++wzKDgRK/5bUCs200abgCaxv+KLPmnlUJQKMLgwUHPvt4gookN6+t
bYYXiuwQxMjmdmxW0JF6uUPku5Z6u8BS/HStBFVHmdEjq4/MhlVX0GKHVX24/1Lq
3c3gZwKsixg1M+lDMK4LfXoRGTzuI80MGJ2RtiQ6CG/QvHbtSy2YQc+uxhtR0NQO
Vegbb3RRY9AQdtNdeWgRe9X6FfYD5b3LdJC03G7tj2BeQIYPUywg7o1AutRCsm34
nIEU02zxEB53Uc/+E65R14wFPga+Ed/g1fEa9JH9imH6u+3hVjqsvbfe6wsRwD4m
jfntOSKuz4YkJQe5/e3cO/VeG+x5EoreoytgNSkbqcEimURYokXvLfQkQYcDawcx
5FeIcLYwoykJctjsmIThMhnS+rq3b8yfmf04DcUfmfLJ1zs78PVdYBP+7cxV0sVv
MKT20tpljUHzeDJqb+/dcshj2OjJSOoKtwP++S/YqAviN8fVsdMgUNf8OsHrxrn1
bQWph3l2g7EYR4pKWSBp+bfSIeE5Aw3M/FeQgpqgjsHxIdwDR1wNn4hXDZb3Mi/z
9Tqgsskk0ppTcFKduvT5RFRqt+o4y9HKUioA4d2oQ8wfmLelX0kpwAWoSE2RLg+p
dA2CPXkn9LNvc1R+kNhwegyeFl8GaDtF/DMNdP+t9703fzQ7vHNj4YbAB1DlzKko
Cph5Eo21Wg9YaJ2cm80AmIPiYymn0sXYvSTHgOYOK4a3AKv9VYpGaIO4RXCv2QWU
CSBIsyeQi8hwaNJu7M9D/1u3PQAg+ZiJw/UgYDPc/6bhL6HCLDRHse2c6p9Ow9/5
8D3AiicCqrDVz/kSjKbD59JBwp4FF0HcGQcU56RU/X1tiTKZSDdJnsFQWd+yA2ay
O9JXsAdddawNq5mv0bL5Wl/X2uPOBW7toK7tpHlY3hfc94w1v/8WmePm7kFIaSuI
IzcITnCAsuXGmCwpaQsmJIA2vBTKidMSTmciKcLGyQU9Qx2oA7zGnMVU4nF+iUEz
HdyJ0eA1fb+L375edWLibEQ9KsWBprQ5oos59CvYQ3gokY9XE90dQlrNtS5oegjO
94SZv52gFhgukGt611CBM1lE89uvQ4AzpXRgw6bt8t0BrHQciz42wVjHLQVv7tU/
lj9zmq73gaCv06yghvVmjFWssm85TAjYxgq7DTWcacsCmCo6pKOVv/H7reDV4qLq
H/rw9EW4WBEp8WVtyAcf3pXjK4W4wAKvgqsok9WxTnpaNm15EOggaKspPCG7E5vu
GVaUp1j5jUXYhXnkG4D/jMyX7rqgpWE9Naz8WuHwjyQvRfqYZWrmBWEDyr8Yz3f4
dBoTi+1dMeqd89ocgProhLZccUrtQdCz8lTBjIgLNVQNMvl33PXeimNRbvZOvqBe
kZadbwkDuHMxKf3xROy1lpyw80Jaf3UL3JPDAub/hTeQCl4TLH6gG46ReFozJrCV
0f6eL6TrYt17+t5EgZeP0cH+ntV9vsUmXgZpEAmtevMfTO4+cuL0xuc3TtSMeANU
0/SQluXUXGMzsEPBW15roI/OAUxIWVkRY/sJGmMTxNTggTAXQprlYJsUN3d3+7BD
a49ROSGMM+tc4W/ewuQFUJc7ShfmM16EWYvt71ZGSTfdhlYwHfIUQIebhlXbEDjy
5XaD0UgYVDePL5gx+SKAtf5W5xdT5VmxtEpmnhTIjyqQtsVX2dF7Jc4yi1ekQ4v+
U5rm9Mi5bHS5KSR733LyQfLr0Ftv2Gb2brvD4HMuzZpA3I8Kn8Kw88r66mEkzAO7
eww3Au4pnVY4INprJVCC4nuzDWZ5JaohfTLc+PXSIksyAtKx2CmjUydjZsZ5Z+1/
4BZ06PDfNVlS17rAZjRUa1jPZzZz2K+IHNEKljOEbj+GlkHSiIBY9iF8CbrjU7ra
WayQiKt4RXYdricXr6XxMR4gx1IZLj7q55wve57JAm8AB7wCk1GyZ4YdgdjCbZpT
f7A34RgZfGjmsnLoW8+OgPh9yQvaoiLRLzqngEFQqELtKmiKVTdcb2CDjE0aYQcu
XsmWtudIkrjuyjFazxPt/veUU3RF7jRYVWg52fvxetmiEuJfRXlITtSbeDgSsx5j
oj/byExZaObnW0YyQbdnlkxGILyAKxF6ZTBrspA3uGefNUhM+4QG88pklSMQAJvE
vcIYG6wlrU/EusUPfk7HdyKLG71EZffMoNHt3tsAghq8sUu0mB5d7d3kpHm7+SpK
g8F++FIWszgnyUc7LPzTOHsEYroRLpHNZ85T2DXDOpsOCfzsZeSsUo7QTvq4DG2p
XhZu99CFzAB21hehTuUyEBwKwgDZQSM1No4AjsGfRxSPAcWwC6ttEmUXPw+ysXhR
iOVYGDkJQRlvT1QVexr0AZowhFgNmrNsRZLMiQsV4yUf6BezVWtpupTCPfIkdm4J
NG4YPHcg/+8S0wly2sf4aUS4t85KfZfbcyRJ8kXRWywGZnq1CdokHZe/nwSCstRt
YPJbcmDZD6rB5jp+HoT4dt/+/J98sfl0T5s4QTV3JpLPbjqb1L/uls4hnaaGqav/
73edIryg9x8DGLhqykL71UuMqdAexP8DHpKt3FWVtzOJad5GbICof2koCSOt7YLb
43Ok0f6tt9kRR8+syhr0ENMZpnXGyYeAFKBLstqRhIrD8xumRf4KVYJvzerhYLL8
R2amumb+d048bW2bS6CctjTH+zv4dhIZMfcbVa8goQDQChx0Rd9v23e1b3tU7jFX
Az2BlywuQRcND9Pmvfx+YliEVZwU5aPZ5d9RNED6jPzMOJkI9Lfk7QP2gUe2cB4p
/vK7qCbnTcGCnqT3r9k+lhPn0j/fiCyJyW+9Ox/WWsXOQrzIOepRZ8+mGf389MHX
DR5R2utJsYF3V238CQ3HUqLvaZXzyl5YihizSvbeGpuo1/uwr0QezZQHdJxWjghc
C9dGp+WSR4WarPiAWKwcOUQ5THP0nbRWqB4vjzm9dek0F0Vyp9pJojJzj8kcCv1+
Qix8NG8uMQBhDJddLimyXXEzjRZ0gmA7MH4JlzGU7YGN2cXZ1a7FL6E6cUpOtSpR
UsdWT2rKBlptlroNMaEMZKJRJuFJwZQZdsfqYfUZGoNkHENS4lpfSL3m40C2ThXe
GQPK3lyc2r9pF3/+dUrncbu9nVFfnSBPndf0T8SlgYX9NVLTFHWLGjJH+xey/Zj8
EuGuW+01m6cM3eocHSXRf1yZUgk6GV6zfTnLGHEy04VXwAcuQy8OtMWnVScvHN36
plt6T6enR3GHHbyqqfDJC1hd3yN874yjDZPjtxOXTZVAcHQGlQPp6hivdyoFTmq6
2k58BJu5xUpa3x3CQBtGSDz5XfDB3Q0iZ3erw8BCkdJsLpAyDlEN28joRpirCwGc
GGZGZeByqbbfVNuJB1oGR3ZgISAbVWV4OdIe9OS0u+VScqhOcin2FmOTO1nqjd2L
3louCmD6dXWtjF2WKkFpwnV4Dz5mUWKMJh5NK+huzAT5FQ8ByH359Xbwcf2gX/YS
0/Fg3Sw5BOGoTijFGByFHFielx4LE8O2Xb9i3peq15NqVbnFonSNYwoB6Ew2zs8F
tBQRK8aG4D14CgXWje8+eNJPi4l7nhQ+k80JRbLuidYJ+GXPNhCm3dBwqEpN1D3R
akfm5naXywo1JKKGCUcFdScXP8ysj3wiXK+ATGaybEl7VukOu6Jx5I/5UVVqOLCN
JC8ZZwb9ouQdZNSjwu9FwmMH/RI96ZIl3M6EIw/rKgcXHpk/TSV+SkzdOY9OiLCh
XKuLXB63Ef9Cp0Lh/VEJktNYrDrT4Vawp/qJKz0cNrZtGP1z16iQ994T0YWdjEqw
ZNttvSvBu5PYsDGmNkV9du+6uRqCmxv4jr2c51r1uFOinoxfnSxS4YJhvMoTq9Wa
EiygwLM0tBUoeklT6RNeJleK7DpgKuYmvpWfGmahlxbAzM6/HjrPp4Hg8ASw+vlq
eIm5CHnaDrTjC6FC90uFfG9bggHhRVoLWYumLgLQpWr/uqkGa5LiYoKt+W3W5rIY
sOu5JMOq9rn1skQY/QckfZS0lQj3lOeBgYhTo0jLP25GJknMpMVg0qvcIL8Uu0Tz
aoMyVqgRx4NFLqBw81hF811yramUwmWN8Q+2rLtUMtn0uGUETXCGtJSkOfbZ9rtM
lR8luwLfjpUYXljxPGeKiWrzRVUXSK2lO2KC3gFrx++D/+ccrOSrur/+oQzUKeul
/HQQxEyL38fE9i7q+UPMn041XuTvtydfWA6d3qHoEP4GkEIHpo9SULsbIaKONwDU
hwzwXwkpFlNnJdAruNDj2/RYWIBRs6TmbDdRhOtqG5oY4wfA6OcteNyp/skTvvSa
70hX7xax22E8Ln0FiZqCyx7aSR1pz/HoMZZ03V/CN6vTqZtaw8GZ6hPHYChN/hvb
b4QnOFLd5GfUH4TltKE619sS7qwurQIfyd+EAjUNKwCmqpRsthgn+NKa5GIDllJI
aBZ6nHobpZL7nFJKx+XPhGUfkwY7uZ1Po+pneuvFKSSvxHUiw17wqN816NSHuM3m
fa6tpju4EBq6affcS7VhmfnSxzB2ew4SqtOZiCydYMSr8AelUgRhcBql1Zsx+ER1
uDY6mGG3pf3bEpulLOYGTtFfn5n3tjMGX28dVaXtbI1XxVmaaP5Jt/l/rAFbbq3u
jgsfRLCIKNsLe9BSpjQnvTAjI4lMIM9hI25Pj9EKCdexQehv9jFCwa4zzLbv8USO
h+ErSzh8kHYk7ulqCGdzvhqQ5JersS3XW0on/gYK12ltp52HfZkQPu3RN9WBgj65
j/XT24ZYqadH1i6QMX4OBic6Weak9SR9ZKyVdIbH7h/Vs+Kfj9Zed+13uv5DLOvv
aFMUitsCKstgzrJJdfFfrrKRD5PH14PvDUZ53xGfwo9FsjcdN8TdqVwSivxBrJZg
5sX6ddVYFbsKUQJIL+RDNihSDwyZbUZv1Esl+wtIvJX97oRUAMID3v0NXFEbvmAg
JhgWqQZjuJ5iG95dOaVF0QEoYNRoMv8GQFeSKikLOYNj8NgKYB9jTZTOVm9sk5ZP
XGAvldGVwGLcuF0MHHLx7XZcIi2ovdrOQ9l4Ar53E+j7GzTOCpYWNjwmJf08fU6N
8/yf+Ons+ijoJVvF6cpCATWKIA0sv7cgjQRRWmu3WLRV2f4k2GDCMM5PU7klwdZs
S0qJsRVNvhujJPAFUQ+bWX4FcTzoYaksPZrjYUB4GWawEGoL6l/ivZW1q1qaZIFs
Nxc3PHYUCp9wAVsArMTdFVWx3XOa88pK47MrHooW83yCQb0ICvdRPb3UHsYg0gGe
vaBhaQT0fubHELPOqq2J8kwJjQTH07Ib9ZKIMMaAtxN7zyU/fJG/XG1S4vLK3F9K
8IZQHZg2/sNFYtBpKMEy5Pt5Ulo/u9ZZh7lzEk3bfnP3qzUSnRnsgUizQKWsd/dm
Vq+/Sj32K3kgnrNXFlXmAkR29yGbj7lADqJaOJnCn9OuOk8eHFd7rU3Ml0b4Vj5g
94XCMG3yFeHl4Z/4eSuxhj0vdIWBCb+IK94lvbTAk8XUaykngHM8A1RU4gkDO3SU
MC1r4N1R3VeD7bo1kVD9GNzpL/mZAAyXP48FPH4mtlq24UCZBW8HFTNd2T7KKqN8
d9MilYIlCDtzpSL6DbAzplzb6UddX0gqDCYT6tr2GWB7iRTA9qAx5JKbdsM7f5S1
pOncB4kH/OLlLRHvoPfcjCvtMuZSwP/GuogS7VumdK/mwgLZA24MTn83wv/4Sp0I
E7sx7bbI20GUoaaNAm1G+XvsHeQ/yYCuJlxV8106OZQyMsGmLuZpXRT91sc0wwTS
qnwl2sOKV3w8LZJKPQaThhD82DgyJsBGWRxALzregnBZ92vD247Y0NleQd7IXW1M
5IrR4k8+OJotZy/9i01fb5KZLUn/gM0XtkY+G/KwrsULX1AW6Y3en79w4YPJsGMY
hnDAqAk/b08U4aKs4Fen3yAQMe+VjiWiUHXlf3h19r9AWIN5Oquo30q6A6ar98xJ
qjP/AHa5ZrflOGWd4JjVHd8/Z85JEa21JIELdv4dOdCcsxf9GCvzx5KjCG0eID8Y
2vGKMqg8NqpJMrb+4GpIGAZHXeqdS4EskRV9eo9mvv6QHKhLer8QDdI1LiD/0YG9
B5fJjleoTWpBYt5ZWI+d0aMc7G2pXcy6dq1jxG3hz1D7Op0i+ftzOQRAFAUfmka+
bXLDRzcM1JUOiDhOWUwIuc85Q/LZ8+IMMQwxdWCN+STEA4R7fDunGMyPonwr+/Fh
CbWh8DYIY+9NWoRLCJJCyUVvKIH1nJ2nnybWN7u1cuKPMIStuq7x2VWOLEmAthwB
wu+NXstpwwMwu8Vw6FG89M3u7XvvP70/q6LpA7rOBenyyx0X2CcZeOMBhW/gjffO
w8cujJl2eFxMpZR7YhlO1sLYefGZZX+WG70l7988zKwK6eQi+Cw1Gx/TTFnGqA5O
+CHTVIpHw2yfaT7ikUlEQ5m+fgjSvVpYfFq38gb7f4+QajVvzDXQzdFb9/T6s9uR
ri2HDsWaVj+O18T9DosjFY2OBpVmdHNrd9EsWQDWkWF3qRc+1PKrSPz1XTwEyXO6
dPUaMsyKPT4+XlQn06ZtlW5aOaDJCcPTaArsPOxH28/iVg48GUdrwbK6r0yrKd4+
pWFbOJ0ScjeSrmGOlNr2g7pV2tLT8FK5AzPst/+73858VzNpJcZlE8/0AFrigflS
/Hyhs4oZGyZ4FLNmv2t2VXXMlpCYADdAgflwZaInbNwQQAw0UJ94atZ05QIEbFbz
i7P+WyFP+GKOYZ5cDKQbUzy0V9NXc+u4gr47hUoJ6SlxQfpLIi+vTLa9Q4NNnQDm
BoQHWFulM8MrLpbvDRzw/H+Uvclsdx7xckPhhhXuWR9DIID0KMBhNfdDIo7I2fQ1
L+uNQwPKwvCszlY45gRva5aCG/EOcXUinWUHHsnPo3cdpxSQqNmmhcuhW8kGUNkS
lIzLqsuy6FhuYQ8Ryg+zem4BaTWsBJcXDUkPB/ZycJHjriNRoERtkfe9RVlQoU8h
IE9aQm0EI6B2uea2pUaroIoAQK6y//bQTEUnZ6tXF0Q6dO79cJMzXSTZ4cwSiGqb
fmIjqV1JiFTzHjupSV9AKJSAiYLNfm32Pw+32v5fxT4zOPtia8g1aAhZOKNreU89
6He6wE0Fv8ljWEmSl/obW024yn9NBkt0kBe9cVuCpjCogb8pTL3X/DcuTeXNgZGS
15rTWCNRdxN4P1JBAacyWHmWX7ET+iCXwEfbUjW2govkdfLgi68IxKSlS3Mep9ch
ecHeZ6pY9VRsWflKN5uXw51nHbCujiHaeje5oetOoGVH4ooCI9UTURQHbrXikxIp
R3cilDIeRPUBiiH1IEGiJmgyMdFCBGQEtiszqjycTlkO4313liIsesZVYzakFjgG
FJpJRobqNzKTdVtHY/bLxByKRwmVrpWZgawCssdPnuui3S+cX9afj8Ge44WKmvR8
QelbkNJakInfC5iaMzDeBXLEz589kCrzw3PW4NlD1lZZeASNXvPCdnYTUKVotHGu
HyVPyqDgYKEPp+QHFoDxmW2ETpfw9D64ArMWnVYVIoqCd+9uCRjQKb9N8AbahMoE
jYlWBH0ptZEfSCEEz/gCrjMrkupz6TwrUVUU7kztOP4bJlQ6cRI8su6+ZoW2wj2l
AqNGzJECDcY/lvoGpC2jl1JA+8s8py0RmREmhanZs68dfsI5SdpnklFW41ErDeAZ
wQUnC7OsWlXFssmNmHyFBpdEXG7J8pvhxz5hEWLo7RUMaBnQLoB47DMuYmTlSKtA
Q6KWrxigDd9KEi+ME6jwE+lkhRtS+JIgmiYbVgJTUeJ4hQ2JW1ztAzoSgINHaak8
bMW4FzE4xwT682QzHvSlLsYxbqA8JJrXKFwD1vLqWU5fAF8icXc/4nvLwMAJI1Vu
kvm0IskG9eJmwqYHKyMzhrP9nPd2mYPDg842HoLAmv/790RclKGIB2afg/7igUx1
Lg2r12MtEFvKo4JrqUH+ooWNTpl/FM13vfkVdQi/MKhW4pfsneYrQnZdy0I6n0ZV
15azRad9XxjpwNDLcrnq3k4uFef/ogT5Tlch0h9I1dkJwV+x3X0j3WjLls7R4UsL
XgxfTVRH2HuIpqhip47e4Kc1K/NhRSaxsOFg6xNJs0mPBSi6UkGtU2+gEv2qU4k7
XBLZw+0blHxWnDgJtf6XkWFf2pkgMnDPt46jFOb+E5Wny47RCm1lWaHNmMvAzPue
NyfEuOEHD3iFBFGw5Ls+qQH1KMeACNadEVw26ZZJ3VgVJdoTQwN/THPMEkN3wjqY
DMJxY2drF59s5kJAwi2KtM8L2M9W3fL6KB9wT7ChERY9UNA6nu+J7CWSz37r1FIt
EeQLSQ6B4Z7Drkrl/qXsv8iha6xMfjZV7rqNE79Gsf3pC3hfc1VxbIcg75dXHDnj
w93zTTyKnwRSUxBBt98aoho5APuWpwDZsXg7VAGBuAV9Yb2XijH/02esXLtrFq6v
1FWhMKhPZQ2/1UsOL4VirgLVHfQ1JwLawbGF1hJVAyVhpsQFSOPikz0cr6DXnrZL
CwtjoiykYu+KsoIT/DcCH7jC490ljVm2ZNv7nIXMOf0mMXojMAyMmywhl1MuBjz5
pJ9FcpTtUg9+SiPFJcN2mpH9/XEfYVbf/BPqxGTU5P60wGeMzT9cjWXUJqXKe+UP
UsbeBF3oKOiy3LVyEpmOuco8KTuqxfgHDlQh5ifm+U/3/SMqqN3JKlzSORfF+rIn
Fy1OVwXhVlzvDOnzBvjkBV9c9HOZRd5gBj5vRDWgZj0bUuVEmfFNgrV2iPl48GGJ
UcEAYxCXzZGT5yR8dRQAXEVwME4m/cHp67lxb2/P0FuLGKXUgPKQaeHDoajrRM+x
kO/0j11afzLW64ZAYB/Wd2eztYYdIUWt4l/1NitDuyPnv2IB6wdfmYmIqx2zbIJy
KQFCXq+yO52gFsmcCmuPLr23Rjqg4mSKPHwegMn/zGGo+a4an9YGw4pS+Cdr43GX
qBNn+brkLgoI2eSvjxTKJ8hlYhJ/7Wwxbdb2Ew6Bmf6YF/JP4wGAo8ILOFvDckPn
X4dXlKNjAxolPZyAv9H/5nrdiDSiVgdr9tkLXrE1zNZ7L3IwVGHC3hLBFyHCmI/t
AD95xYdlfkL7CL20L9h1YoqRPKGOwy+UOHWOi6M7S8Oq4BE+L7G8t/RhjOyq+Vcr
bAWhKv9qO1d3dm9y+Z2PR/RS2bt8M58XksdP35ekD5rUSYLXRSINVls/GOPwI0aw
gXJLzmcIeCue+reoYWboq9mhofNdlpG3Zpd7D3x7sCo9iSExb6B//1RpqkLSMavH
LwIkXx2JJTsWmdjBPt0b2Tcm46O5SzXGAx8DRB3Bg+lFLVscBlta7aBqEQJUfLMv
QRk79GpqUO6OzNwdmMxn7RZtw4i2DM1huc8ZO4T95u9K9qg3a758G4D8k7FGpjwu
lCxhL1siu4PYNvxWWqE6j+NYzEdtjiNKzKCk24Z9xztujmhnFSb12wxwaIpbabRT
ccC8/IWAnK4FCCtBU7RyIVBiPiC2gjaMwfrdEVs3ruLajTFbmU7oKidjuQcVaAjT
IZqs7bg2Bn785XZ0V8UAqR6CLq2/3QnEyICME3DdJvgjthcHp/6LLQcww/cSDN2w
kDa8UWxEbjVaOxwMmzRbrRpWJGF90FpKNen3JjLFOZ/BbXfpntbviZtAHsN6bKUa
JnNuTQfwXy2BnP92/QetDLrKf0yND4iIXrp81Ondu1Vhv7v33K4a1kbBthnL/BdU
+x+JExrAkUYY8B1gW/B+R+fTAkuTKUJu/vZpWYsreelSggqRiuJp2o/vU9+8XKid
OrW6ldlrElD4LJYeo8u75p0r91lLu3dYv2NBrEFY5B1ZuEZEU0EybcWbUpt2ftdc
Au4VUd549bgVgGkFKVn0rylRyrAdHiyPBZji55sXiMCBbDjprXtPsJtdRICfsaJE
2HwcNX9bokhKPu0CzEfcEfvCwJZYvNFGJWMVs1Bh7eVKI3tNci/SHH7OL0kb5O8H
185vm4o67eCmokoRJryLH00/NbBttsVK4COhMOAvwXAHTbwr397OftpCP/EGJkQp
eCPlyIq0LUXrKggmcULkmQ2DSDIfbP7SX62Xb1w2qIUMWYnzvz4r/JEis+ymdbeV
W13cv6rBgBkXGrlIsfdhK2U/b3R9xonqZddMNvSAUloQ5svXfF/s3vMvZw+Tzcvg
6ZFSfqyiKu5nUhBdo5G36KgXk3HQMmqB/wdQtjsTA+ChSp1i8oCc817W5xpo3Ztm
fKKV3x9b6/bQb4hgS9xCyPsjvKbul/B4J6xDhI1qTPK/vVRQNIJDGpzp4PxeYPVx
kcjtbqjVUt6nWTq4LqYEmKZ6ob2GSH9Bk2uGGzTDSshL/lQecxNxUCl+pCOSjzNb
g7gQG05WQ5aBi7CMhYYi04b8NdVBrZ7GxGlfeWbvMY2OfYZ2QsYuAzeAlDbtSa2d
rZndEgM9d/0Vyr4vVe11UAdqXejkiF5OuLu6pn/cGjUEf4JA4OJH+v5/WNqYELd9
nJpkV4cXmd4I5z6fj8hkYK0vGdAc4Vd325fL+MjLjWxuaG8jpOOcou2jaZ5Zj2J2
sWqp71CB3OOZl/CqwLFCvgKNTawOfqu2XsRAZaZdl3su1LbymR7sWTfP5A+JTJFQ
JBS3SjaiGZc59uwQfgsytcjnaRdEKyhiBtqy/H1DP+AcR4UZ6RZugW48chPC4wrx
LKOFua+0/IBMd66pTAdaCZ7ZwE7CYDBoyFlfutsVM5khw2XrFKsh6AYiJqxGX+yB
eqdaXt6ivb2RQ7ct8S7tk6Bg5dRMeOJF9VBURDzV/swK4wJ29PxDhDHfrkcHKlim
qtbHkwEPTgfD3ato/tSCTNTV3jxXlpfKQ6k+In+FCngj+hxrYCz+MKaTNE+gxxQM
lWzutbsgAp+LyGNZkQRu6b847SY5ABuGUvrBLc5oEAOfSJeqLFNB9l5iewJ3Bgii
72oSkhK4NpCpYBTwo/2qhOSY5l/ozniFqoE06ItM4uDCOjaC1yeyCf2YL5rKADdh
d/ARRbP7CWzgrK0Uehu9VDBdWbsGdpBweK0YQAUT4ADo8553HG53o/Hs7kjbGadd
UBVKYyTgGSlARfxF9/ZlvpeK/y9olwjuHgbN+9gT0aOxGq/j0nXL+kQq9KXKet+n
vXTMUFtCjMXcVDGAtMAEh7Iwf64D7Z46pzDDJ89Py5S2BPKDndAMCakzCnDqBzt2
moNW4GD5Wj9tNSiAcSfId71oKr0MViF50u3Y6ablrKIrlsdiEQ7ZY+cKJA3zAeCW
QyPIkYAYPriYm3ZXA4o5AfJKySNdP0OlTB0joRqNG7zRib/gt46INfpb3m7Bf/XQ
kx0RcxkHEW7KIU8g9e6B29fWj8WrvrqeQjM30Ut3ElGq9Vgmgy+9SmRaU23B1o7J
WeVLO3nDOL0mFkcEGoILUwhJFmf0JSMkyCnaUb0nPd5rJJpZK9I0MRM2Y9VB4NiT
q0eW8b78FR0pkh5o6Oc4w5JvR6ecQe8cVwobO5i/M2O4Yqgp5xcNlCvVRP8ilWDW
MGaeVg8zlkZoxbdcFUbyQjrof90XciKDapBGVaT7Q2vRXJ6Xo1cID1d9ya1ETBCy
nqIPdD30WO2jGuppcoHmZpnKUvdxhMYcD/uwr7k+zz1Ulf9ETSXLw9DtBKGjAQxf
EXFOE90r3SEKWVUIBB54OqExhb2lYNJ1pdZ+X9N1BCUC6M8MIMOZJ2ZzH4QEwAjO
mBx2sWMdmSe3n0hBU/eGTO8FNiVXquTqDc7ydM0bfxM6sHO0SXAtGrgv/lZqXOlX
ArAVTRSl6vcmCJqsS577J+H/45ULdPx7BS2rSzHGJj6S+8nD2xtJAgWvUyXq3CSI
eu64NY+CU8lAFbQ7xn8PWRaWC5cLqlN34kpdPpJQgwf4Yi0/13wURLqa6BpMJpTL
ehKBa/kQj3qzq2JtRhclvRI5KZ4eqOW3g1ulDGZwUQAkGjbsHeHcjJIzmLK/j8RU
5vyCaNqBHXwjwQLJGK7226fQq4IpYejfILg9vUm7i6sC3punTEef5m8jnaZrzyDP
6ok5C11C/Wr2QPieiZWsoDC7E2LJbOkd5TYfiYAYYcKp5AL0Izem7vYy6CY7jwIF
tJHIUnNTM4NMkiXsB+5e/dp+2bsHgXSPyM1pPPHgJjw1PuM/ze1U8EVtH1AKg5wP
xSxGOt7Gaqr49e45x7EkUCRtlaQsCGRphYcE1FfWpmKhYVL5uX5vUGDme+dtndIg
nwNR1KqMNXtNOXlMD0zbr7K+PjMWtO7p66NtNv9chTq8jKPJnj02LZ//cWO9AXFj
vWmuB5iQyVnpglp3Sgc6AXN8kgfX6wk2smzKNm1qj9+o7lCTxXUMwdcTXZWktU8u
iY/ERriOxbsaB0X+i8fmSu/H4cMN9OlYKWVIDRzZKHVcwpwgsbWxBQaQc1buwn43
busBbb7zJE9YfuJG49pO69eG1tw1IQoJFbq9EyjuHZH7ryoK3hofpgaVegUmnt88
PYz6K7AfGqs0UygQZRWFmuO5+UjRxdXvPuA+7ATzqohkK6sGHmIxTus+QbmV5GzR
bvmtSJFT5W6bZl97YMrKLO7jcxZWKLQn0GU8V0yAbHEwUISxs3ajGYRoTXroy3E1
6YW4aA5Wj1wiRc1AjWrjZNQMk3Ix5PCStMldTPJjQcFZolc94jto5zBT0lA+A3Mh
5XDHJDPSGuL1riz+OR1rcSfNV7RcNdZ3GA5ewyF2/RaBg+GowXdvFseOk/VoYsdV
ksP2GNp3m9y24twH73dKaQBvGp4e+v33Um43uCyZaebgK8gB+4di7MtzSq0FFGT6
7RKeXAgNjgCH+8tX+Jr5+vLaiFg/LMjOFaZqrGAMbpfeJDS4koUr8bGzhwiuwNeu
FI2GJlZf6JV7Qm3Xj3zvKdLH0LWNlH7EJ/BVcQQ7hCgqsdI4FPw/TtcVNZGRIiei
KmNqZOWJKgqQ4UutoITw0a1Tx9HNeauQuA+UI7Qtp96mIKHqEh5Qare71T1u+V5A
RUTbdGFEHuH9ZDnCu2hO5HODiZG6ZdCaowiZN+LALiur8xu2JKR7Qcg4P3eb/2jw
QhX8tdWgjga2kzodAY9WNbE0xlyXpJMI/foXiGcL5t0EwcIu6+7ki5Q1xB2xQ828
K1Tcs+Vy/HpHJTyxH00o4ufmzi0hAySCyxToaMycAgdzxRnlMDMqnFLUcQ28yTEh
oMiKbaCjJrU46M9FfY4RPKQlKu1NmQjrNCsUKwJxUMLgR+HSfGanA/E18dd+it+h
XT7uHLoe5peV1xgK7ywV5xLxSxqtE3qJxd5zrW9CQBdcrHDd1dxCvdEWV+mZfw+x
SM6shsy3FcsO8gFTQE9HTOqkIO3mgB9z40xwFoamtmQA3Tr29xIgALb5Or9iElW7
YhnGUeR7Lkg2JBUUxTOJCrqQ5VWV4WyF+EilsEfiU0e3hEcqvBfNejAQWE1bAot0
FsNsdnFn8SxYJXTwHBPdsktK0bKACwvEuYYsoKNTua2uq/w2iElhOoixn48EtToR
QJgWJWGsge42uq2xafh2TY5F8ZIio+dt24EBg07P+0dPlKuQYe6cW4JfTFpqleSv
rXhrKsQFzCfP7dOG7OUNoBCQYe6IEy1yAbz37V455+lTCgqwJaF7X7anIYn0kZXn
/wfj77tiubNnml94B++IGv4gjjJk4Qmy7dfb4Pf9XOKFjQbqJ1Lp1aZ+LqAqZugp
lN/FN3f70ap3+Auu1H6lPHePq71vq0JGLtqBwsFL9q+NifvngDRpr+Z/Htpb8kDj
7xGhuMBiyFKxT5x1MdBups1CJGLkEzM22JKH2PThIZRGhgPCtORx9FRxJY59NBXO
5FCwhu95MrqR0YyXkyFwwEeAlnSX+PLc5UHBbhO7hbvD/JWums97wXrTpSDZ8KKM
7vwHaKWvTSlzWhFE3g5npDbkFCjwfltlbXG/rRDsNhd6swa/JzwjCXsKuZ/7ydNW
e5eoX3PqBbRIov0b7dBN7rs2tgJqkkVD12V3GIPxbOk/dVXSgyz/Tfo4XZE+kOA7
KG+NORiVbQxhp/GZh1s4GJ2vbGzpOQ9h4bcUExwyyzGqq3x6hiDYytAg3XR5W2za
NzoquVdLFLD58L9PT1YvgrAqyk/SkC5+Ql1udzXDYGvEXGyrG8pCNel2dVpgFxQ3
pQklX14cVpl5BTavclGqNNkq5LlWpGIPt+4VLNVAEEkmWWfgolAYI8yL2SkZ5TTT
Wu1i/0NiDyS0SKfpYAVqfrtPS7GvZ0/dmFAR55qyb0XiweJnOqJgxpG+EnaF8zqf
XOohNdLHmvLHmSXRYzoEr2M7SIOg/EXxsd4TXckri3IK497ylYtsj2bdnOYbD1MZ
11TsYyezU5q/rtoX4Dgl2P605zN3vae7HeioX5bxByZab7gMFe9MkklMiWW2XE8y
U3MvDUklAoRBu7AFsIPmDAiOIItblA8eSQj5aHba7V3LOC1pD3YtEFVxz3lScnI4
twq2T/BjFIl0VHsLKYRFAaHR7eANZ17HJrzd+Uc+hWaJNRf6IFs5CTBkoVzaGVmB
xRRl8uB9Yim3cWpTO2VUKctBLm2mjrdywtxga1H5iDgUSiW7skn5AXoNbvUhECWc
O2Rclcf1X35j6mutufRc9tXu0D6K2QYR1asshroGESUFtop//RHH6oJW3G05kypU
mo4/qc8+DKtcQtJBtnVhJFwB1wQOKjCwK5bdNNU2JOY3aWZh5hTnltofTTylMmot
CdS17/1XVHNSNtTGscF8MGLd0HjEnkIsjQzONcTfvXze+MZ0lT8Lnuvwg0oUXwCA
SJiBQ4wyGcMXjZw1WE74xkQ55svnVd7xg+nLlRgs6H45MhYYHaYvehpl1rEOnC+Y
c5HQCFTPgfHkcw/RgVmOccy2BG9FhwunZLbbr/c3NiHATaLRa0Ibg0Z9x16eHSin
PDKHKfRN3PNVKDyIdjZyANhtW8IAhhIMPJtX4KkLNOgukxWf4rD0qim81Wiak2cM
kRQJooCPiWeQI8vJ6zNxKKROXV/K+tHazdd+/RDRdpHdU6HdxFYlkV0bUsrQmO+9
SSnl0k8dUSwwMJbqZIFVjhSwp+S+KQgM5v5aSya5UzEBjW8GosmDNghOp0m+yzTm
nKDXEHFNqWE8iij2VD0KpkwHhD0yapHc3MYCTKH/d9FIC71hVSb6AyTiLQfHZ0Ib
LKBAphyzv6aUtgVLY/1tA78K5f+f9q6EIGhWmkqQKFzJ7zgd717wutpsdC3kkJX5
JRstx4CJfFPVOHAtf+kRaLAkVTQFl9u84m/UOlv2zquKBy7MkhCn04C58gODLtXX
4P4bqnRpwIbAMTj2P3oiHwVinVZTn6rR+FtmnZ915Naqs94CG4Dq2qu3WQiOF+G0
+mCmxYDBzfAzTdXsegDKSsdtv6ML5j4TH36L/JbPrw0wRx+T0EiR9aEzoHlq/5uD
AVioDofUzbLNlFuzNVBkAjd7yLxYzL9SSwczaTieHUR98ZfYIz8DjVmfzdPK5iCb
SFG1Uoo/gLS/ZG4fsNGpOyTkW7I99nnTppGcLvO5N5pLbn78kiSqfNVnRIcDp0VD
YG8KUaLbYi8I/0QTAUxJ50WnlnLzqz0UTB86U3YZ0LSdHsHvmZuaE0+BscPQ7Yym
VapMtpU+AtRsqu0hWNdW4hFe5UPV/RPGDDQiqFVv7VUbiMbnEEGeEllL4cRYQ5K0
ilRN0fRXnmZYFlGrKXaLl/jF7iuidWswFG/nbvpUQAIdn0d91qcK4HNx/z2QZvp8
RL7M54J8qL9Iswn1+SpTXkStByR4YOtzYWCFy5my3rnTEEUgIra9DjOHpVVZQSXQ
TUbWj+d8S6VY85UeLhJJDW3pMPk2qEA9ooG8VN33B1T4ot0UbuK9tknhoLhNpwMh
Mzx5XXwLY1whVTMUnED4HpWElLi+1MHt9LFdlmYMCD48aQB9dQ1gVQLU6R8975JS
0J3BgDkhUcIu2LZtFwZeTRlLrZi7e0wn2NoHa02zcMxNI6gnCESJdy5J+khEol+D
ZREOk1J6pMXSEe247v85Miyuv/A1+6fgyPJCtJNWj6z+z7WQoSVDE/PMfcI0z6DA
F4Ei4YhQztYZxh4q7ctbvN0u/YvGz+0i/EAplSw96kBTs2K2FGXgR7dvlXbtnltb
zNE5OgOnNocaWTF2Wiwn64b3awlaQuFT/WvYF5xbWWfXwz6O3Ye00ENBLB3C+etF
OF9ojQqD0bcAzJN6t9yMH0WoORmeEE3kj2uYuKjx1ag7nKLMGrkw4oZxEXD1elke
KkS0awdMLEooE+dGgcK/EgeX+qAZfC1UlI+f0lAMqSxUP40Hey02STGLnbhohebQ
xLU5QjBNqrpm2PT0UW9TB5MwprCDgFQWMXGz4WpqzApBsvjJE/iNDNNaSoZSnksM
GO3WEkEQ+hfjBy9AjJByxKSA/4F7xP5b3aOf1C9GpboxDN96/40T5AJHkOOk1h1x
anT/KdAp0CSW41i9wq0wsyhx8gLHwnZJameVlcklyzV0ELOCW37ZdOM1q14e+Hsn
dTZ2YzFvlrEvfcA5empo1SYuVUc3a0j5sM0Vzaw3oWFGbgj5rh8weu8orYNKvg8c
aI5jaOqQGWwra7Gcb9lBGhBNWOnhLNJBWiLmhPDfG65I0lGu/TX/Za7AqmXGgPt5
p9D2/cM5JAv7Uqs7axtrPwg/OO3tZWv5ldjclCv4uBNOTgBjLGlKcf/RodIcV5bd
baMC1aOzT2lrhy72M1daTRETmos8Tz96kGRweE9RV9fy5K7SalLSZbgHjQmdc5rZ
JkxVt39+TLBd+EmPpgiJ8MnVsxte4D8prrT7Q0e0PwoRQfcvzA9wwQRzqXdsdHMV
5NBw63dlSUJEQhLYWU85PD5rJIUSPrCsItE7KQ2CDQ1nYfS1qRgK6mK1TBumvuwh
SlZuB2ykXhh68dDoEL2yqzS2rukQdRkNad3oI5/+xDPAMjUWcCQ5S6ujmTkbCdDq
6/GnpsITek92FI0xXO1jpQh55VRrtziEBBjvwyLVFvx+ggsd4W5NSybFPJiicTEv
2IVWHxd7lQjLatYEgQRqNNKPcpg+ny40zU4vsLqKex7CAtKG434QUgyBnrdmwu71
CrEtlDCdgnJR0ztsKrT0a2eazH8chXeIGsnPIci/pqWFBmRsXEsBCRPpkYIlOLG7
e0Qn2NgsaE15LUfOCXCRUoT50tLtB0d+CrcLweMha3AXfkPi/XhoBDt9/RP93gcI
SNANoYRb+B8uIgpWnGOIbeoxeJX5Lb2F+VEGygXoSb6E7Eyu6Ltge5RDtEeMeNiD
zgxtlyQ0ve/Z8McAbi802Lz1bo9B46blP3LWojcC2a0ookZeHs4Y1cYx9gyW59dl
xHeFBHpnZieC6JWWRghOTRBbKd0j7Ew3OksuOvCBffrymSoSPgDcQud/1qCG5Q9/
FjXwIaBjND+UIbPGP8kAB6Q96pO8HJENIc5qJcl4v7bRmhQEi5yKRrTH2fYo6I78
ckk5YBpyjx3pYpXSM22dUCvkMSKsCktK4iHE8gGSKidakGS8LwDXPo+esiI6YQ4r
DjcFzVvvuPpk2wwU1qV3VL8kIQ6+3ohGBdqUmhfA7lwMgQzHpxcfw16seP5KkdPt
NDn5prcmTBai+QAQV7jQ9G8rYtSX0jEpGMcK69KaoQtDA4Aj0oSAkYjHpNgzb4W0
/3BBuL0Xii54CdRh1y/jH04Sj/b/1qfx6V6JOULEt5T5BvdoYKb+AtFE4qLcqj2f
ceg5RXj96xkRNvU0XmaoZzAJuHqzV64G+ZIZkn6gBFHZhpzq6h3rVUiRS6EAGtYO
20kCVPEQP4lQGfl0g3vbpiipWFA5yuBh4MiBanDMdU66Qjm2mw1TzOzlX3lSZSL8
3SxHeJaesLZorEeGvQHpik7tax47KymzBSkRq01XyfcxJj0c5FZtfqHxjE41W/TH
bzlG7VXTG05De4QSSC6hI1q3AecxSiiGa7HpQVuCSZ/RusTPEcSXfH59eHhK6Ft9
B13LvdNrCeIVamN99sPjA+Ci/kv4oIRfEkYu0P1wg2JmslVq75Sz1pC+YvTPXlfE
qYaJ406Hf203J3iTtm2hoxuYa7GbIBcCbh6NOjZ1UKjpp+swQloxLsvigqKww5VB
6DWJkuWt4F9tS2w+hyBPJa+nfV5+N1eZUsgknl0EU6OLwsJAyZwupZLnl+67Sb2+
xXokQUNBIHOLyGAZV9k198Xg3X+0Cef5GzSrLh3+6qsxh4jcLrtScKIcKZV/ZK3f
jmxutOfWJzyt8k2uOVT4qitT42b1MjDKsUlZUJZM5y7EviYjHZA/l3MAWf6obqiI
H7h85bha44EIrgBytd7ks8NamEe0EyZ2uOAAwPRx+POnGjyh3oSA6YFhK7lHitjx
pxB+K+rvv8RO24qJmpEYKgtWYqGR2GDdZWNuCYXm0SvEZYwGcomFyFbftGRmCpzs
ukT0nrjg5Lp9PXHQsdK1GHV+IDLIQOf1C+Uv5oztOwGetl4h7ScqRSZngEl8I/og
bd+mWpKw9OlCHJ7Cf1gV/85ejfZt9WwAw9uFDcpCaBxavUUxSIIho33Qu+oXAu+v
MWL4kmOxza9M1pabrQxSeXM4uq4ebh4VUUiQ7PjJPGqqyEAGwjbPzPrDZYTzJ1z3
wtvEQPm5w5jvhj+3A7w7KKX3WTWgWr3y1R8AXamqiSrwHGJhtooPucw0YfRyfp3i
vdEOywOD5Fc0Z/GwZOpnwienINopdHBdUl20mKYIP7gt/OuDd5xMR7jg8p8OQZty
veIW4mfhBpK/HR3MzQRQvbF9GWOZPvZuTDwKlt5+cuz45enxdtwZKwTApiaQCfHs
h1IC7njEtPpFuAStgPxjCPj+TomP2gsNUZXVy/S/dGYaXGT06FZSFFkWEgfyhj5j
yOWI5MSNV8J7gCVnedtbf2w1F2lrecNA1QnzCJPIz/1keVnz/bA20dxEv9UkbhpL
ZC2VydCUO96aa+K8eUv1Sj/HJyRHtcyjK1vSXZsAbaWLDz0/pb15Bpwkn1Wb8niC
8rd34o65J99eEJg/TDelVF7VfonKPHtpLVMF8MfNSNTciNuaXgAM1Gdoow1JTtFY
T6PsC1KNOyaTv0AUd5aDBdmE+OJPzJJ079zE3gY06NPhohZly4Czwb1XZyApDQcm
QOXNojd1Ul8f435H0Yd6ROsIzSV7U6SXBkmuuYdnxztGzhtmTK7X+zo6L2dXJuGb
eb0YgexnCtVG2VqDrWOGakJgEYk1TuTCKsNyHPqE5KrC+XvjJhLuusPso2zsdEmL
N0f4cVFqmMgy+qQOPX3r7ouBbFWq/iBiFA8zFaZnew2p2hvVCAP5WwifLjEQkphJ
vuw89dnOGAWTO572V1A1lAV5q1cbWvFlZDtuMAIGZ2/uN+/RlojHcwOnixE29u4k
KNaWx6euAhD7htmmI6nHDiPLulld5ZHehGtXbD8NRwTlx8yE7/pq/F1uG+gFCQyS
gSukHE+Vnfaex0UOVTUxiEHTpoS3U90X+wL/aMlAneWQx/ObPtc3/uS1WjxzF8/5
Q2N7QWwZnGMX96VpL6CHCX9TU2mythfTLz4tM9LsbtyMJ/8/p8xTMRyT/Madvd8F
u0DdxdgEd0qGxUI+DzFwlxfLNPFs7US+LkkaxjSqpq0CB3mGs7h/gG/NoFtzwIfq
lt4oTj7HEV8IeP61bMkdJGnbzgo9hfaJnDQfj75nLu6fPpFXdQmhaY4NH08LkwrW
dCHxnMMlVIz37o9INoPeDPziJ2BP9Ut/hQDJhEhlWu6bKvZVWdh2i0pt9/6DV1YS
lCM2fi/pou94pqT9kIM05IXDgjqq/+9yE3rVqUYvaQ4pZZvUVB7PZDChHEmMX9NX
fBNEOxo81LTmaus657jwtcMiA2jX+ntkLUR6gu9i7kVGieCWXpiYEcHx+yunUUwN
1OfZFEBj7RFEDfMuRB0GhiO4R/EG9e2OqpG1oWwsfIUYB/pMLLLsnxDaj0wfVmeT
PXXbby243QPke23GiyF8N85iEQ3Cfm1QpzpIkKOUqb/xq+VzlNwa/I886SvXA8Pm
f+rEnSzHR/GjqBZZS3Vy2kT7zUxb+ajj1cqPAqJhQxPqH7AUL4yGcdCmZqML5Kt4
HN6LjuQTYfMj+QcoxCrQ3iH9D8vU5VU6Bcz7se6f/8BtC2dDcTFi2wM9AFX19G4+
BpQy7UgLh2sw5P2jh/cUMUL24vreRimlWOV1ClwELDHZ77Ojabn0a4v65tShdql6
gz2dcrsvWRGfs4ha9gNo+XSb5+hpQ0VeMRCj44gapCCNWDd0xCMvdd111vEzge7j
U2ryLLycgA5wTqtsJK4AbuTxfGcM6JM/5oOSVQ/eCZ7xl0Ah1hBeS8724psqvQMh
yzgLZyDXVSz4LjYKhqDIjH18CV8fuDZaT8PL0z8S17VRFn9N4u5Zq7+iGtzLiePn
Yz7c0zvWfL/y1PdkzrwZv/aHTm9iT5eIlvar+IClzw5oulbCSIqbjMK7tDbZDqk/
7nPSmNTn5Em9m/amKysvJv4hQbKppN5Fi4z6dXC9LEiB2OOyog0Agu5JD1LU6218
jCFl6LKUmXQCPlIwhVLf+qPmHC4322roEFW6vj1yJrDM9/6TlNovLth4hQ6ZbGPv
B65wCkSrMyY5EmibcfCrfqzsv1HvTjIibvoMlGXt6FclpKnFplgVjQIoKE02bkGA
NOCDAX7Vs8FTN1RdKxzyWZ6xpADkbv+bz4wu7B5D6fDnyIUVAChpKggNa0ohnYIi
0B/j2BpTMAwH7duuvRSHzfCMG1UiSb5J3C9fA/EYiZlGWk/dl4Xa/9SNgB7NuqHu
gA3Ruf7rK14j3YVDPVJSKl6KgGXBDuyZOwFJOjpx//3g+iETt81G0rkfcP0UnIzM
Y1iQGo8gjtGxTb8zS3R6Mz9GdUCcf0MA0QBtb3u6IyPk9ITppRogumx6Vh2b685y
N3hAipH44SSvoDZ5T77HfiCTF1VQE3tHgijQ08nC47IHQO+TqZzqO5V+mVGvfQf+
XdxRLhzRCFvGHBlABRKkfJR3TGSKsbiQzNjUDXG+PDbKwcKm43pFq3xHaVkOv70/
fh6n/fanZyOC3jBHFh0jjLQwhyMUbgCaY1TH2fKo3PDZLnvWyuZpjy8vkD+zxZE1
oKuLHwYu3h+CWMj8okG8R0vs5cppvBI0iHvcwIpgEbpGO50rTBrQtD1vKn3UA1m2
uCe6FIPyPnG14hmFR07edM7S+YJxpl4X7EyOvbv4iD/ZU3dx0dX2BbM2HRPOKoX7
K31bfg7Mn8Uo+8b1J/7qT+AcPcHRAunHJzjgMzqY234Maza0r7TanxW0Oy8/sQhO
maV9BHbF4LnJ+uhkRPzFTyeWyJYpIigzCWhU6zNXVD39TnW2rjpULcB54gFB1fCr
Q16gJLkWZaI/kOOSoshg86kbfLcdypLCsPa+OaK6Xp1M3FwUPeWd3afSUUgzaVdI
C+OlpnH8xV4X5HIq03MG9+udWS6tbABKyVIcwKJARIGhmZ1Pg6+LiCPjrcjGfCxj
hQ/Arxf+HYrUhIn1H7zQDWK+IqaVv/w/s0MEw9uAuNT/pTcFeBDrpIvricN4lDnr
aCHc6YXB/XvAlsEEi/G27mT9BkjZGmOaITcgSEkegSg67qhaRXer1/csPgyv97lC
845yU/h624U1hgKN/oHG2NzghOsgDgEpmB02aQAn2XcFHywQFiGIezVCDIx5BlWk
dtTCDteHOsaoy238Q1fdNudneEg3xUuNmc4qHiwyYUfP11IDm5VGkVwCFIGHolKz
7Rwr+hDHmSG9qJCzgb5ZYCWQFkqtEfWaw2hI8mZF5W3yRSxZlB9Arm8C2V9xLyB6
6KZfcNPFJvN0Wz0SuVKXlnLPsLQ5H5HWyJriiqW0ay0TNXL52uJq+tWr4LfqG3Tp
5ix1DYSmMVh2i32A98rfscET9Sg1Gjp/iwerGnsRixIciehG850WwdUgbXB/uNp0
NcIoMOWFEV9ih4PfOBgJnHtym+JkOQ1R4WCrh24DOR8+kMOVWMSJqayO+ObHPyjg
UEhuwlWqXG4oS4FBtVd3kbw8a/l3fT6PR8JjsNgY8pseI6ezf15y5QsRomRBpSS4
RWQziuMRNYBdIAyj3tNPSu9VQ1OY8Hu5r5sIrfJCgMC/MJyK2O4b2gG0e4fqeRBb
Bbflmqzq7NAVEQptbliikcQVPGSQdv+Tsez4tYxw53MKLakPAVjtzdcU0ar9kDdS
mIID6AR7I+gdGAXjDFsJsZFJxgpgyU0ASxDilwkmOc5wBic6xVtNlyLoBybt3bH8
8JEC4btCnKVX3YPzt9h27EuXAcM3kWp4UZWefs1zDhqSLfmI2rzQFWBZYoQU92Qu
h7tJcCm1vwELfSNIn7QVne88xWzej7p4Qpv5qB6lZyqsYr9LTH0nRkx/RDuXmRE9
igPr34dbm55q9J7eLl7z3ls0b29kxO45oTb5/RrV0/Sd9wRaPBkLhITium3Vhc39
c87hCJqBIhfTE3zdFgdYI0UPRXP0rZbCMsudTYq+5iZTelabSmEJLT9pYFDBYPyu
DR2kXwOJeipVO9wJCBvoQiN00FjZFqXDdXXpknG8G41Xy4KJr4jEIj/aIlLwI1Tw
cviUkfUhQHr/QYEPV2eRl+ZKDqLy6cyiuvo/XVwR2g13eDz/UthgvJI0lT9nUKyy
HKt06lM4J+wMpQBLM0WWYWvwlFheU29YpduLYAGcWtUPE66LCg8IdBxTWKmlTPHF
h/3FDs1UgF9gUW7PwbtZV/lnlHiQJeg91BvK1/KnCubEMhaEb2nUCUk2xky6atiS
kO/ot8arJIE1c+BMyg56UYl+CSnyHg6u9KCFpd9q6ARbAY0lggkTvILWRlnmQrQk
GggrTfjooBl8BImWijJAg5Cc2x92BxD8nrCPJghxcRgY7b8t4CgF5qfaxzwDNVpP
0gDR8DC52BAC74AqdjNdu0sPv13BEPzMmhwkCFvqYW/HQeL49n6sZLGzf/4H1drF
phtZKJ11KlFxbjChzdjovgWLA8rhHJ/+EdmnsN1VvFocniRQgDVAJCRPVVh9bP7r
ZOS6l67nwP4dcCOvRKVRe7TIbFkaYp7iB3jhvb9W2IvUD+nTxaMn1yK0X/LJtlcp
B0Q1jCizXfvqCDuO6K2QMtieKcEJW81718XOYOkX7UqpUwXxdiFb+G+U/zHyzAIh
fiWOcX1cRVF170QQMzKy/MKGXu4Dxch6es2k9U9u0VxikTvJxQxo+1ZLalYgF6m8
AkgigMvMnekfZeZGEeph4yNOBpZNQWpMImwah5IL04bdKcCovktnwKHngPA5IJm5
nqPhAETus3gj63ssakWbKprALTE7tz4ZAYhmjpmLSEACI0WNTvoP7dE6qLUUsgih
tsi3Yro7Ea4/3gponMSjU5qAHQvT4EvzNTb68MVsUgg1Ua8z+Cz8DV9A6VZznjio
ICk1/J+SvPdLBi5VKauLLiHhzsVWy7nLJxyKeUs/ne49gSwzHK3xht5rzI3svXja
tT86aHlEQfUvZoxtl2PCMfz8IoZnN8g7hZIUEKG4kS78HjrZXMywdh4NN+FgcKxH
CC29UvQJ+TblfYgMCrkNqi+TymkVHMdv+zkXf+B0uRBYpgvaF7lxVUuR6FS9zG7u
c6mBNBO3/+5wT3XXjn76DbTkOsVpQxk6ytTtDcLOb+irsyE9T+H6tPoCDn8PHBFr
ojHQCJqhvRJLItOgLxds+SbSDk77ru6APV5Pv9AE4wlaaswrj3tMhU42i1yFgr1Q
6VaofqDYKlES2dqtwM6zociaWx4muqZXBekWF52PBny/Phau+j1jwj6kz/mIVI8/
Xx+VI2dQxk1yCTw/GUVGMqeWYWOsYM6SkQiQG+WtZIFBZZhsMbsKFuj0k6vaU87I
I2daN2pXNfB4f1kcrwk9dl1qyFD8peCrbW/zjPsN7Vc1N9uzFCvKWqNv8Oi0ne/h
68hg3apEPmCzn33/d4QLEmR5f2s5rVk49QqjZ56HslKTDaFV87hDAVlz+5fBaNYv
HUNcIfpb/WozKriIDXTejAbWBDZrB4TyGFSd2kn5AZ2ZN/nDY4jrNsrZPG+Zxek8
gE5dLhb6asoArVvMT5pCzngOidIAqiPbqAcmVIEKhcmo7zzIA+mp50VTKibEnbp4
KM67nnKIXfo7+gagV5V+YNZWW9+RVG+Xn9XsDYTTNYHCc7JHWsxZkkOSN8k76ovt
SenHSreLSdhHl9k4nt7Ex2oAZD8hN97ch2adPs1X5W/GDTGSMoctQDcjYinNa55X
JRspMZbeGQOpNclpZk4ysb0ExpIxNFaKtJYpMVPdkIHzFIgXWS+HyIDOEEwF4Qi4
sGOIsr6ZJMZVsBmLh6P/jD/4GFGUoBblOqBLcz25oB7mpeOIxqozGsJWcH6ZzBV9
cdW0rJ0i1PZaQgriVaS4VOXc1ufM3yQCooL5PKZM1qNvMPUBZM5RFvtS1YA/09zC
jIlOPy3+4J0GIzn5JIrUpBvh3kyOWMpU/8V1+j2z876xV9q+/EKaJSbwcAHCy/a9
HG6O03/jVCQZYA3Bq0OAAThM/G7drF0LkU7c9FoHM/NDe7EtO1eIPq1hVV3ScR5T
vzXMGRnsze0r9LD81M2PanmBOGF8HOYi3pTL59mHe9LY9D1Ix6fKNyS3ohgUtvLu
C8Ne14FyA9HSGyghOOejDZlEPGM+vBZMwzpQvQrOUwqJ2VSMZNpxy102iTcGXGIg
Ne3bC001FbTFIvtdkJ6iy3MF2EeN0dUA0B6fi/GIpjgeJ54PzOGXGEMPohtNe5DK
+4Uuv3AquDFhMhN/DXgB4CXcErggnklOG5NzJxrAZgamrk+Zt1pEtEhBHeboA1vW
cwszRJRZA1IwrEcysMvlx5B2W7l0cweNMJwXum3ti0/EDURmxkqFwZKXoL9AZ9Oh
NOsqa52xNmpS0OSQxfiFHyVNoPVVmEqX6l/lwMDrVcKnbSOqfd80sFrbz40qe94m
aspQ7JCk0izpCIsplnPABA7m5xtyWXYlIy1s6j6z7jyFWSSJIAs733U7AMuXJT/n
PNG9EKJmVXtXFCx/VulpeVLKcVmOa/JZXh7KKovXDhbdTTMTN/qkJG4uZ/uo0TYP
CVyNmlQCrFPFt2LZz73RI4jHUY75pEKw9BrPtJnZCHgt+kQ7P4PyDO/TapsPuJFQ
4FU8NsBt4j6mgQ1dxBIEH4TAAr5oIyzMTKdQnFlZGg40smiphl6tu67sWSvBtmOT
rLc9Ius9bvk1nKy9QOT40OmNdvoA0lVjuHOkNtXxc7PtmV6rDneSypsolJ3ioWWS
iemWww3U87AlLrKgC5PP7tD5TuFbtF+7ZWKxWD61rHBdffvCstFvuZfyjfh61u/K
mefDhxUasqjnjQFO9Ct/2YP6GUYNx6L/+oqJOlWo39CEkhgB/MnhvGEgMZck/EK6
XbOWut2D3Kkl90vxtZbMNIzuO6jcLqTwzzTiNc5jMpC//p3ktz3MsVfCDfz/VlBV
0Kdxg2piNKSBZhZ4OKXYEqsyw2xJjMeFL2v3SZ0k0q5+mcH3f+9ma6Z28dEIeX42
DqQOTbW2+pxcKA+MnWiscDAVQ6JZnqt9H/2bXlkbTyD6byrTNAzwGZDM+BYLnYqU
p4n9f7jNEY5ZCuVnhbTxLNIfQG5gt1bS0G5FhhohUJLQzCXTsaQTniWMILwcx9Vc
oYAYUmexc69xz33fXphspT80xiItZcsz5PoJt6a/mWLxAmZsrPD9dfzuaYT9dEBB
k6ck8ZGkD6mtsH/f7bP3cV4RdlNNl0lAwbpzbNiHjGvn69n6zGM9T13UhSmqlH3c
AtIuw9z8QSXKOyoOTPys63DzoV9hI3eI0R4AzpqmCe+DMCs2IGfjgrXdeI+S6zQg
WmWOXpCONW76JrVKTQ+y4/RfOeAJv00E4yDclGJgAdcTafCIHL3sTvtljr5Z4k8C
SxUAKF30eqiHbTaKESBqEQYdD91Ffv/JQ/vIQDLymptelvIcaY1ZCXIg1Xk9szDO
/+PrxRgHoNDSbEf8SNGfKzJLO5Xzh9JwBo1V/4PbEzKDkFikyogFzHscdVhWcMc5
k6gpBkIXDHXPOao1166DwjH0XYL0Pbm0qofiuv620j9xGpjwAw1X8qsvJiP0XZNN
7KGj0jQecYCuoafpI8DL7r+AqPzs1oG9fbQXY29du2AL0RCfLbLs6xAmX+mT6cuk
koJ6VdM6YWSREn+oZbneYdnhdU6a04R8BFc5/WtVfSjrjfz2UsiKJju6yAVepQsd
x0DEp4dM6HAjqjK1c9wo2UDgef6h7J+kmJs/pdxGX3njpLsa0zuf7QIPikVUmeyx
CKMaFjdsKVODt7o7xjs1nvN3hd7Pm1+jJreJLYss//DKifi4vAphmCoPfA2fw8Uq
4Gq7iWWU0lRP6f6vPVMemnggYuU8UyCZK59j2e6PXZ5nWv2EVBMTaSb9W64Hh9Bd
3PC/QU5pwn31yF2O3zlSfOw5puYdbVRNXShFUAnR8q2BHBDDL7o6anK4gbkDauw+
3yIqyLMO04teS4OidyTWxgak+yBn0W85IL0zdzarsKP/jiQ6ZTTAia7/wsgD5nWu
+o2XBIuxyZQpFhr7S1+c4q9f/M72r4qgmYIfJ10WvyTOXi/w4XQZUZZbWZiPfGrI
p70FqrqZDYkTczMfasPN55SCdM171M6HpuUrZOTs/GlYs9ysboStFQYvd03lIeW6
kegJR3cuM0F59wXnO10mcP3SUlVkVwquJo7dGTAjnUcZteUVpB9Yz0Rz1b4cEmrY
FJm19W3eagGVGD+E92z2EM2bg7KV1FZGUjvQLsjyp0vZsNHJEDbsXuz+IsCZ5IpW
HzSnFChV8A1kuiEq0G3Oaafr6S4r1JwnhO/SFo0RPxVnCdAdhitnTVr1P+gVxTgd
CGyqiG+ljhQWtYQ0bVkYL6eNGJt+gOb00Xfa9KblH4FQg1f3Q68zPbdA2nVK4U3Y
FuX2MX3VCwessYIFYqxRHnGO0xKwfc4t+97ROmnEtUgnsXW8BieZhiIZOuUAJnUs
y2/ndfyck2RwnStxr+jImz4oOk5Y8TWm+Nq0hgCrsyk0uEjCC9UzH5Iiy562lLOX
cBKtRk0D/8LTzCKIl7u4DlkgZ/uSuYrUcBCSfkaszI2EFEA6dWWSFRelLEciRcet
chPKyCZPJjMAvsVWuGd7BF8D/m38VhXMeANgvBNzyJWevFfxIc8R+UpDkebkNkAW
mObvlDiWXTiIVNybmDni4RMD/6fpprSB83Jg/xQSbyj6HVyI0w2YPM+NlG5XL/Yi
R2yhNh9kerfBlDWbvF2hRpIRovzdC7Vzc1YYhjhQRtXEyjNAZVXNC5/3sXyovg/s
D5NsvW83kTZU9mSO2c+gwpXhV8MPiBz42/noNmybPTH4iU3jhqO8RENghBGbN5zL
lTQdvTlJG6sQ8Kx1C0AnHUJUK5sEiuP754iF9zcu5b98JNf0YmL07O7nnuUXrryz
MQUCwH5cMWNk8AL5ssGH5XwBBgxtQ+h8H5xmTvXSjZQ7vpRfEuVCmgLMjMmwJlov
1hDRCipkOX1tSNcQtsU91WatjxCesJpw2JK2bVFDaqBDSqw5ueDQG2XWYmmQhLyb
nnqJmSIjWetjtn9XwSeOtx6OhmkvJ55/1QGwhPNvBXIYq8CKCSKoTFjEytzq+fuk
BJFpQ1tsgqbs2Dwg6q3qRCN1KhFVuopetKg/+bi806E5xd0lhZjzub4/ng3YAQKZ
MhUxHyVIsgbpM0J3lX2zHmE9ny0fMhez/y2n3JT48qc=
`pragma protect end_protected
